//--------------------------- BASE PARAMETERS --------------------------

`define     DEVICE_XP2

`define     DEVICE_FAMILY        "XP2"

`define     USE_HARDMAC
`define     NUM_POINTS           2048
`define     MODE_FORWARD
`define     SFACT_RS111
`define     DIN_WIDTH            16
`define     DATA_WIDTH           16
`define     DOUT_WIDTH           16
`define     DATA_WIDTH2          32
`define     TWID_WIDTH           16
`define     TWID_WIDTH2          32
`define     ADDER_PIPELINE       0
`define     TRUNCATE


//-------------------------- DERIVED PARAMETERS ------------------------

`define     NUM_POINTS_2048
`define     NBY4                 512
`define     SFACT_WIDTH          22
`define     LOG2_N               11
`define     LOG2_NBY2            10
`define     LOG2_NBY4            9
`define     NUM_STAGES           11
`define     STAGE_WIDTH          4
`define     NFFT_WIDTH           4
`define     WR_LATENCY           9
`define     HMAC_NON36
`define     BE_PL_DEPTH           3
`define     OUTVALID_SEL

// FFTC2048_beh_all.v generated by Lattice IP Model Creator version 1
// created on Fri Oct 22 10:11:48 CST 2010
// Copyright(c) 2007 Lattice Semiconductor Corporation. All rights reserved
// obfuscator_exe unlicensed version 1.20aug2009
// top
`ifdef HP_FFT
                                                                                          
`timescale 1 ns / 100 ps
module ls1e5c2_FFTC2048 (
            clk,       
            rstn,      
            vkb84a0,   
            rtc2502,   
            mt12817,     
            hd940bd,    
            tja05ef,    
            sj2f7f,    
            qv17bfc,    
            lsbdfe5, 
            qgeff2b,    
            yx7f959,    
            pffcacc,       
            wwe5667,       
            ou2b339,  
            cm599c8,  
            encce40, 
            os67205,  
            an39028,
            fnc8144,      
            vv40a26, 
            qi5137,       
            bn289b8,     
            en44dc6       
            );
parameter pdyn_points    = 0;
parameter plog2_points   = 4;
parameter twb8d6f    = 0;
parameter enc6b7b   = 16;
parameter hq35bdc   = 3;
parameter hqadee3     = 1;
parameter ptwid_widthr   = 16;
parameter xj7b8d4   = 4;
parameter rounding_method= 1;
parameter pfe3535      = 0;
parameter gq1a9ae     = 0;
parameter med4d71 = "ECP";
parameter phard_mac      = 1;
parameter pscale_reg     = 0;
parameter ptrunc_laststgs= 0;
parameter vv7105c   = 0;
localparam ks882e6 = 2*enc6b7b;
localparam ngb984  = enc6b7b+1;
localparam vve6110 = 2*ptwid_widthr;
localparam db84433= 1;
localparam bn2219e = (pfe3535==3)?2:((pfe3535==0)?pfe3535:(3-pfe3535));
localparam zxf60e7 = (enc6b7b>18 && ptwid_widthr>18) ? 5 : (enc6b7b>18 || ptwid_widthr>18) ? 4 : 3;
localparam fc3fcb5 = med4d71=="ECP3" ? (phard_mac==1 ? zxf60e7 : 3) : 3;
input                        clk;
input                        rstn;
input                        vkb84a0;
input                        rtc2502;
input  [plog2_points-1:0]    mt12817;
input                        hd940bd;
input                        sj2f7f;
input                        qgeff2b;
input                        encce40;
input                        ou2b339;
input                        cm599c8;
input                        lsbdfe5;
input  [ks882e6-1:0]    yx7f959;
input  [ks882e6-1:0]    pffcacc;
input  [vve6110-1:0]    wwe5667;
output                       fnc8144;
output                       an39028;
output                       vv40a26;
output                       qi5137;
output                       os67205;
output                       tja05ef;
output                       qv17bfc;
output [xj7b8d4-1:0]    bn289b8;
output [ks882e6-1:0]    en44dc6;
reg    [ks882e6-1:0]    en44dc6;
reg    [ks882e6-1:0]    ks3b5bf;
reg    [ks882e6-1:0]    mrd6fcb;
reg    [ks882e6-1:0]    phbf2ea;
reg    [ks882e6-1:0]    uicbabe;
wire   [xj7b8d4-1:0]    bn289b8;
wire   [ptwid_widthr-1:0]    wlbe0cb;
wire   [ptwid_widthr-1:0]    zm832e8;
wire   [enc6b7b-1:0]    iccba1f;
wire   [enc6b7b-1:0]    yxe87c3;
wire                         ic43e1d;
wire   [enc6b7b-1:0]    gbf8740;
wire   [enc6b7b-1:0]    cb1d024;
reg    [enc6b7b-1:0]    nr4092d;
reg    [enc6b7b-1:0]    sw24b7b;
wire   [enc6b7b-1:0]    hd2dec2;
wire   [enc6b7b-1:0]    xj7b0b4;
reg    [enc6b7b-1:0]    dzc2d3f;
reg    [enc6b7b-1:0]    wlb4ff7;
wire   [enc6b7b-1:0]    xy3fdeb;
wire   [enc6b7b-1:0]    shf7ad2;
wire   [enc6b7b-1:0]    dmeb4a2;
wire   [enc6b7b-1:0]    bld2896;
wire   [enc6b7b-1:0]    pua25bf;
wire   [enc6b7b-1:0]    zm96fd5;
wire   [enc6b7b-1:0]    phbf55a;
wire   [enc6b7b-1:0]    xwd56b8;
reg    [enc6b7b-1:0]    vv5ae1c;
reg    [enc6b7b-1:0]    xyb873e;
reg    [enc6b7b-1:0]    zz1cf94;
reg    [enc6b7b-1:0]    qi3e535;
wire   [ngb984-1:0]     xl94d4c;
wire   [ngb984-1:0]     xy35331;
wire   [ngb984-1:0]     ui4cc50;
wire   [ngb984-1:0]     qi3140a;
wire   [ngb984-1:0]     vv50285;
wire   [ngb984-1:0]     iea17e;
wire   [ngb984-1:0]     mt85f8e;
wire   [ngb984-1:0]     dz7e3ab;
wire   [ngb984:0]       tj8eafb;
wire   [ngb984:0]       qvabef4;
wire   [ngb984:0]       fafbd2e;
wire   [ngb984:0]       psf4b91;
wire   [enc6b7b-1:0]    co2e45e;
wire   [enc6b7b-1:0]    hd91781;
wire   [enc6b7b-1:0]    cz5e07e;
wire   [enc6b7b-1:0]    rv81fa0;
wire   [enc6b7b-1:0]    jp7e838;
wire   [enc6b7b-1:0]    dba0e32;
wire   [ks882e6-1:0]    fp38cb5;
wire   [enc6b7b-1:0]    bn32d7d;
wire   [enc6b7b-1:0]    tjb5f73;
wire   [ks882e6-1:0]    go7dcff;
reg    [ks882e6-1:0]    tu73fca;
wire   [ks882e6-1:0]    kqff295;
reg   [ks882e6-1:0]     neca54e;
wire   [hq35bdc-1:0]    ir9539b;
wire   [hq35bdc-1:0]    gb4e6e8;
wire   [hq35bdc-1:0]    tj9ba2b;
wire                         pfdd15f;
wire                         ipe8aff;
wire   [plog2_points-1:0]    uk2bfe6;
wire                         fn5ff31;
wire                         eaff98f;
wire                         ldfcc78;
wire                         the63c7;
wire                         mg31e3e;
wire                         wl8f1f1;
reg                          vv40a26;
reg                          zxc7c69;
reg                          an39028;
wire                         vif1a71;
reg                          ou8d38b;
                                                                                          
                                                                     
                                                                        
            always @(negedge rstn or posedge clk) begin         if (rstn==1'b0) begin            vv5ae1c <= 'b0;            xyb873e <= 'b0;            zz1cf94 <= 'b0;            qi3e535 <= 'b0;            ou8d38b     <= 1'b0;         end         else begin            vv5ae1c <= xy3fdeb;            xyb873e <= shf7ad2;            zz1cf94 <= dmeb4a2;            qi3e535 <= bld2896;            ou8d38b     <= ipe8aff;         end      end
      generate         if ((twb8d6f==(plog2_points-2))&&(pdyn_points==1)) begin            assign pua25bf = xy3fdeb;            assign zm96fd5 = shf7ad2;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end         else if (twb8d6f==(plog2_points-1)) begin            assign pua25bf = xy3fdeb;            assign zm96fd5 = shf7ad2;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end         else if (pscale_reg==1) begin            assign pua25bf = vv5ae1c;            assign zm96fd5 = xyb873e;            assign phbf55a = zz1cf94;            assign xwd56b8 = qi3e535;         end         else begin            assign pua25bf = xy3fdeb;            assign zm96fd5 = shf7ad2;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end      endgenerate
            generate         if (pdyn_points==1) begin            if ((twb8d6f%2==0)&&(twb8d6f!=0)&&(hqadee3==2)) begin                assign fn5ff31 = (hd940bd &(~qgeff2b)) | (vkb84a0 & qgeff2b) ;               assign eaff98f = (sj2f7f &(~qgeff2b)) | (rtc2502 & qgeff2b) ;               always @(negedge rstn or posedge clk) begin                  if (rstn==1'b0) begin                     dzc2d3f <= 'b0;                     wlb4ff7 <= 'b0;                  end                  else begin                     dzc2d3f <= qgeff2b ? yx7f959[ks882e6-1:enc6b7b] : hd2dec2;                     wlb4ff7 <= qgeff2b ? yx7f959[enc6b7b-1:0] : xj7b0b4;                  end               end               assign xy3fdeb = dzc2d3f;               assign shf7ad2 = wlb4ff7;            end            else if ((twb8d6f%2==0)&&(twb8d6f!=0)&&(hqadee3==1)) begin                assign fn5ff31 = (hd940bd &(~qgeff2b)) | (vkb84a0 & qgeff2b) ;               assign eaff98f = (sj2f7f &(~qgeff2b)) | (rtc2502 & qgeff2b) ;               always @(negedge rstn or posedge clk) begin                  if (rstn==1'b0) begin                     dzc2d3f <= 'b0;                     wlb4ff7 <= 'b0;                  end                  else begin                                                               dzc2d3f <= qgeff2b ? {yx7f959[ks882e6-1],yx7f959[ks882e6-1:enc6b7b+1]} : hd2dec2;                     wlb4ff7 <= qgeff2b ? {yx7f959[enc6b7b-1],yx7f959[enc6b7b-1:1]} : xj7b0b4;                  end               end               assign xy3fdeb = dzc2d3f;               assign shf7ad2 = wlb4ff7;            end            else if (twb8d6f%2==1) begin                assign fn5ff31 = hd940bd  ;               assign eaff98f = sj2f7f  ;               assign xy3fdeb = hd2dec2;               assign shf7ad2 = xj7b0b4;            end            else begin               assign fn5ff31 = hd940bd  ;               assign eaff98f = sj2f7f  ;               assign xy3fdeb = hd2dec2;               assign shf7ad2 = xj7b0b4;            end         end         else if ((twb8d6f%2==0)&&(twb8d6f!=0)) begin             assign fn5ff31 = hd940bd  ;            assign eaff98f = sj2f7f  ;            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  dzc2d3f <= 'b0;                  wlb4ff7 <= 'b0;               end               else begin                  dzc2d3f <= hd2dec2;                  wlb4ff7 <= xj7b0b4;               end            end            assign xy3fdeb = dzc2d3f;            assign shf7ad2 = wlb4ff7;         end         else begin            assign fn5ff31 = hd940bd  ;            assign eaff98f = sj2f7f  ;            assign xy3fdeb = hd2dec2;            assign shf7ad2 = xj7b0b4;         end      endgenerate
      generate         if ((pdyn_points==1)&&(twb8d6f<(plog2_points-2))) begin            assign gb4e6e8= lsbdfe5 ? {1'b0,uk2bfe6[hq35bdc-2:0]} : uk2bfe6[hq35bdc-1:0];         end         else if ((pdyn_points==0)&&(twb8d6f<(plog2_points-2))) begin            assign gb4e6e8= uk2bfe6;         end      endgenerate
         assign fnc8144     = pfdd15f;
         assign iccba1f = pffcacc[ks882e6-1:enc6b7b];      assign yxe87c3 = pffcacc[enc6b7b-1:0];
         assign wlbe0cb = wwe5667[vve6110-1:ptwid_widthr];      assign zm832e8 = wwe5667[ptwid_widthr-1:0];
         generate            if ((twb8d6f%2==0)&&(twb8d6f!=0))             osf5e4e_FFTC2048 # (               .hqadee3(hqadee3),               .pdin_widthr(enc6b7b),               .xj71cad(ptwid_widthr),               .plog2_points      (plog2_points),               .xyadfc4(enc6b7b),               .phard_mac(phard_mac),               .device_family(med4d71)               )            ks15b47 (               .clk(clk),                         .rstn(rstn),                       .ph38443(iccba1f),                 .ri110f7(yxe87c3),                 .wlbe0cb(wlbe0cb),                   .zm832e8(zm832e8),                   .hbd80ed(hd2dec2),                 .ph3b7a(xj7b0b4)                  );         else if (twb8d6f%2==1) begin             assign gbf8740 = ic43e1d ? yxe87c3 : iccba1f;            assign cb1d024 = ic43e1d ? -iccba1f : yxe87c3;            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  nr4092d <= 'b0;                  sw24b7b <= 'b0;               end               else begin                  nr4092d <= gbf8740;                  sw24b7b <= cb1d024;               end            end             assign hd2dec2 = nr4092d;             assign xj7b0b4 = sw24b7b;
         end         else begin             assign hd2dec2 = iccba1f;             assign xj7b0b4 = yxe87c3;         end      endgenerate
         assign xl94d4c = {dmeb4a2[enc6b7b-1],dmeb4a2};      assign xy35331 = {bld2896[enc6b7b-1],bld2896};      assign ui4cc50 = {xy3fdeb[enc6b7b-1],xy3fdeb};      assign qi3140a = {shf7ad2[enc6b7b-1],shf7ad2};
         assign vv50285 = xl94d4c + ui4cc50;      assign iea17e = xy35331 + qi3140a;      assign mt85f8e = xl94d4c - ui4cc50;      assign dz7e3ab = xy35331 - qi3140a;
                  generate         if ((twb8d6f%2==0)&&(twb8d6f!=0)&&(hqadee3==1)) begin          pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           shfd9c8 (            .clk               (clk),            .rstn              (rstn),            .din               (vv50285),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (ldfcc78),            .dout              (co2e45e)            );
         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           ec824c5 (            .clk               (clk),            .rstn              (rstn),            .din               (iea17e),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (the63c7),            .dout              (hd91781)            );
         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           wl80422 (            .clk               (clk),            .rstn              (rstn),            .din               (mt85f8e),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (mg31e3e),            .dout              (cz5e07e)            );
         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           aab9f03 (            .clk               (clk),            .rstn              (rstn),            .din               (dz7e3ab),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (wl8f1f1),            .dout              (rv81fa0)            );
         end         else begin         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           rg5843d (            .clk               (clk),            .rstn              (rstn),            .din               (vv50285),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (ldfcc78),            .dout              (co2e45e)            );
         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           fc1b64c (            .clk               (clk),            .rstn              (rstn),            .din               (iea17e),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (the63c7),            .dout              (hd91781)            );         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           ofc692e (            .clk               (clk),            .rstn              (rstn),            .din               (mt85f8e),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (mg31e3e),            .dout              (cz5e07e)            );
         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984),            .epaba5f       (enc6b7b),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           mta4b11 (            .clk               (clk),            .rstn              (rstn),            .din               (dz7e3ab),            .cz709f8             (),            .qgeff2b            (qgeff2b),            .except            (wl8f1f1),            .dout              (rv81fa0)            );
         end      endgenerate
         assign jp7e838 = ipe8aff ? co2e45e : phbf55a;      assign dba0e32 = ipe8aff ? hd91781 : xwd56b8;      assign bn32d7d = ipe8aff ? cz5e07e : pua25bf;      assign tjb5f73 = ipe8aff ? rv81fa0 : zm96fd5;      assign fp38cb5 = {jp7e838,dba0e32};
         assign kqff295 = {bn32d7d,tjb5f73};
      assign dmeb4a2 = go7dcff[ks882e6-1:enc6b7b];      assign bld2896 = go7dcff[enc6b7b-1:0];
      generate      begin         if (twb8d6f==(plog2_points-1)) begin            assign go7dcff = neca54e;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-2))) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0)                  ks3b5bf <= 'b0;               else                  ks3b5bf <= neca54e;            end            assign go7dcff = lsbdfe5 ? neca54e : ks3b5bf;             end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==1)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  ks3b5bf  <= 'b0;                  mrd6fcb <= 'b0;                  phbf2ea <= 'b0;                  uicbabe <= 'b0;                  tu73fca  <= 'b0;               end               else begin                  ks3b5bf  <= neca54e;                  mrd6fcb <= ks3b5bf;                  phbf2ea <= mrd6fcb;                  uicbabe <= phbf2ea;                  tu73fca  <= lsbdfe5 ? kqff295 : ks3b5bf;               end            end            assign go7dcff = tu73fca;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==0)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  ks3b5bf  <= 'b0;                  mrd6fcb <= 'b0;                  phbf2ea <= 'b0;                  uicbabe <= 'b0;                  tu73fca  <= 'b0;               end               else begin                  ks3b5bf  <= neca54e;                  mrd6fcb <= ks3b5bf;                  phbf2ea <= mrd6fcb;                  uicbabe <= phbf2ea;                  tu73fca  <= lsbdfe5 ? neca54e : mrd6fcb;               end            end            assign go7dcff = tu73fca;         end         else if ((pdyn_points==0)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==1)) begin            assign go7dcff = neca54e;         end         else if ((pdyn_points==0)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==0)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0)                  ks3b5bf <= 'b0;               else                  ks3b5bf <= neca54e;            end            assign go7dcff = ks3b5bf;         end         else begin            me5334a_FFTC2048 #(               .ba99a50(ks882e6),               .ho69416(hq35bdc),               .gq1a9ae(gq1a9ae),               .med4d71(med4d71)               )           qv9fe30 (               .clk(clk),                        .rstn(rstn),                      .pfdd15f(pfdd15f),                    .uk2bfe6(gb4e6e8),                 .neca54e(neca54e),                  .tj9ba2b(tj9ba2b),                    .go7dcff(go7dcff)                 );         end      end      endgenerate
         ea78733_FFTC2048 #(         .pdyn_points  (pdyn_points),         .plog2_points (plog2_points),         .twb8d6f  (twb8d6f),         .yz26d41  (hq35bdc),         .xlb506c  (xj7b8d4),         .ip41b33 (bn2219e),         .pscale_reg   (pscale_reg),         .fc3fcb5(fc3fcb5),         .gq1a9ae(gq1a9ae)         )      rg5282c (            .clk(clk),                     .rstn(rstn),                   .mt12817    (mt12817),             .lsbdfe5(lsbdfe5),            .hd940bd(fn5ff31),              .tja05ef(tja05ef),               .sj2f7f(eaff98f),              .qv17bfc(qv17bfc),               .os67205(os67205),            .qi5137(qi5137),                     .ipe8aff(ipe8aff),                   .ic43e1d(ic43e1d),               .pfdd15f(pfdd15f),                 .uk2bfe6(uk2bfe6),                 .tj9ba2b(tj9ba2b),                 .bn289b8(bn289b8)                  );
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            en44dc6 <= 'b0;            neca54e <= 'b0;         end         else begin            en44dc6 <= fp38cb5;            neca54e <= kqff295;         end      end
      generate         if (twb8d6f==(plog2_points-1)) begin            assign vif1a71 = fn5ff31;         end         else  begin            assign vif1a71 = encce40;         end      endgenerate      generate         if ((pdyn_points==1)&&(vv7105c==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  an39028 <= 1'b1;               end               else begin                                    if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                     an39028 <= ~an39028;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  zxc7c69 <= 1'b0;               end               else begin                                                      if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                     zxc7c69 <= 1'b0;                                    else if (ou8d38b)                     zxc7c69 <= zxc7c69 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                                                      if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                     vv40a26 <= 1'b0;                  else if (an39028==ou2b339)                     vv40a26 <= zxc7c69;               end            end
         end         else if ((pdyn_points==0)&&(vv7105c==1)) begin
                     always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  an39028 <= 1'b1;               end               else begin                  if (vif1a71)                     an39028 <= ~an39028;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  zxc7c69 <= 1'b0;               end               else begin                  if (vif1a71)                     zxc7c69 <= 1'b0;                                    else if (ou8d38b)                     zxc7c69 <= zxc7c69 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                  if (vif1a71)                     vv40a26 <= 1'b0;                  else if (an39028==ou2b339)                     vv40a26 <= zxc7c69;               end            end
         end         else begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                  if (vif1a71)                     vv40a26 <= 1'b0;                                    else if (ou8d38b)                     vv40a26 <= vv40a26 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end        end     endgenerate
   endmodule                                                                                             
`timescale 1 ns / 100 ps
module me68523_FFTC2048 (
            clk,       
            rstn,      
            vkb84a0,   
            rtc2502,   
            mt12817,     
            hd940bd,    
            tja05ef,    
            sj2f7f,    
            aaacedc,    
            qv17bfc,    
            lsbdfe5, 
            qgeff2b,    
            yx7f959,    
            pffcacc,       
            wwe5667,       
            ou2b339,  
            cm599c8,  
            encce40, 
            os67205,  
            an39028,
            fnc8144,      
            vv40a26, 
            qi5137,       
            bn289b8,     
            en44dc6       
            );
parameter pdyn_points    = 0;
parameter plog2_points   = 10;
parameter twb8d6f    = 0;
parameter enc6b7b   = 16;
parameter hq35bdc   = 3;
parameter hqadee3     = 1;
parameter ptwid_widthr   = 16;
parameter xj7b8d4   = 4;
parameter rounding_method= 1;
parameter pfe3535      = 0;
parameter gq1a9ae     = 0;
parameter med4d71 = "ECP";
parameter phard_mac      = 1;
parameter xyadfc4  = 16;
parameter pscale_reg     = 0;
parameter ptrunc_laststgs= 0;
parameter vv7105c   = 0;
localparam ks882e6 = 2*enc6b7b;
localparam ngb984  = enc6b7b+1;
localparam vve6110 = 2*ptwid_widthr;
localparam db84433= 1;
localparam wje829b= 2*ngb984;
localparam bn2219e = (pfe3535==3)?2:((pfe3535==0)?pfe3535:(3-pfe3535));
localparam pf611f7 = xyadfc4+plog2_points;
localparam ie3efea = (xyadfc4==enc6b7b)?enc6b7b:pf611f7;
localparam zxf60e7 = (ie3efea>18 && ptwid_widthr>18) ? 5 : (ie3efea>18 || ptwid_widthr>18) ? 4 : 3;
localparam fc3fcb5 = med4d71=="ECP3" ? (phard_mac==1 ? zxf60e7 : 3) : 3;
input                        clk;
input                        rstn;
input                        vkb84a0;
input                        rtc2502;
input  [plog2_points-1:0]    mt12817;
input                        hd940bd;
input                        sj2f7f;
input                        qgeff2b;
input                        encce40;
input                        ou2b339;
input                        cm599c8;
input                        lsbdfe5;
input  [ks882e6-1:0]    yx7f959;
input  [ks882e6-1:0]    pffcacc;
input  [vve6110-1:0]    wwe5667;
input  [1:0]                 aaacedc;
output                       fnc8144;
output                       an39028;
output                       vv40a26;
output                       qi5137;
output                       os67205;
output                       tja05ef;
output                       qv17bfc;
output [xj7b8d4-1:0]    bn289b8;
output [wje829b-1:0]   en44dc6;
reg    [ngb984-1:0]     fcb8586;
reg    [ngb984-1:0]     zz16196;
reg    [ngb984-1:0]     ba865b7;
reg    [ngb984-1:0]     pu96dde;
reg    [wje829b-1:0]   en44dc6;
reg    [wje829b-1:0]   ks3b5bf;
reg    [wje829b-1:0]   mrd6fcb;
reg    [wje829b-1:0]   phbf2ea;
reg    [wje829b-1:0]   uicbabe;
wire   [xj7b8d4-1:0]    bn289b8;
wire   [ptwid_widthr-1:0]    wlbe0cb;
wire   [ptwid_widthr-1:0]    zm832e8;
wire   [enc6b7b-1:0]    iccba1f;
wire   [enc6b7b-1:0]    yxe87c3;
wire                         ic43e1d;
wire   [enc6b7b-1:0]    gbf8740;
wire   [enc6b7b-1:0]    cb1d024;
reg    [enc6b7b-1:0]    nr4092d;
reg    [enc6b7b-1:0]    sw24b7b;
wire   [enc6b7b-1:0]    hd2dec2;
wire   [enc6b7b-1:0]    xj7b0b4;
reg    [enc6b7b-1:0]    dzc2d3f;
reg    [enc6b7b-1:0]    wlb4ff7;
wire   [enc6b7b-1:0]    xy3fdeb;
wire   [enc6b7b-1:0]    shf7ad2;
wire   [ngb984-1:0]     dmeb4a2;
wire   [ngb984-1:0]     bld2896;
wire   [ngb984-1:0]     jp4f44a;
wire   [ngb984-1:0]     med12bd;
wire   [ngb984-1:0]     phbf55a;
wire   [ngb984-1:0]     xwd56b8;
reg    [ngb984-1:0]     jp4acd7;
reg    [ngb984-1:0]     swb35f0;
reg    [ngb984-1:0]     zz1cf94;
reg    [ngb984-1:0]     qi3e535;
wire   [ngb984-1:0]     xl94d4c;
wire   [ngb984-1:0]     xy35331;
wire   [ngb984-1:0]     ui4cc50;
wire   [ngb984-1:0]     qi3140a;
wire   [ngb984-1:0]     vv50285;
wire   [ngb984-1:0]     iea17e;
wire   [ngb984-1:0]     mt85f8e;
wire   [ngb984-1:0]     dz7e3ab;
wire   [ngb984:0]       tj8eafb;
wire   [ngb984:0]       qvabef4;
wire   [ngb984:0]       fafbd2e;
wire   [ngb984:0]       psf4b91;
wire   [ngb984-1:0]     co2e45e;
wire   [ngb984-1:0]     hd91781;
wire   [ngb984-1:0]     cz5e07e;
wire   [ngb984-1:0]     rv81fa0;
wire   [ngb984-1:0]     jp7e838;
wire   [ngb984-1:0]     dba0e32;
wire   [wje829b-1:0]   fp38cb5;
wire   [ngb984-1:0]     bn32d7d;
wire   [ngb984-1:0]     tjb5f73;
wire   [wje829b-1:0]   go7dcff;
reg    [wje829b-1:0]   tu73fca;
wire   [wje829b-1:0]   kqff295;
reg    [wje829b-1:0]   neca54e;
wire   [hq35bdc-1:0]    ir9539b;
wire   [hq35bdc-1:0]    gb4e6e8;
wire   [hq35bdc-1:0]    tj9ba2b;
wire                         pfdd15f;
wire                         ipe8aff;
wire   [plog2_points-1:0]    uk2bfe6;
wire                         fn5ff31;
wire                         eaff98f;
reg	[1:0]	bl5f6cf;
wire	[1:0]	vifb67e;
wire                         ldfcc78;
wire                         the63c7;
wire                         mg31e3e;
wire                         wl8f1f1;
reg                          vv40a26;
reg                          zxc7c69;
reg                          an39028;
wire                         vif1a71;
reg                          ou8d38b;
reg   [ngb984:0]        wjf81ef;
reg   [ngb984:0]        ir7be3;
reg   [ngb984:0]        wwef8e7;
reg   [ngb984:0]        ble39ca;
                                                                                          
                                                                                       
                                                                        
                  always @(negedge rstn or posedge clk) begin         if (rstn==1'b0) begin            jp4acd7 <= 'b0;            swb35f0 <= 'b0;            zz1cf94 <= 'b0;            qi3e535 <= 'b0;            ou8d38b     <= 1'b0;            wjf81ef <= 'b0;            ir7be3 <= 'b0;            wwef8e7 <= 'b0;            ble39ca <= 'b0;
         end         else begin            jp4acd7 <= ui4cc50;            swb35f0 <= qi3140a;            zz1cf94 <= dmeb4a2;            qi3e535 <= bld2896;            ou8d38b     <= ipe8aff;            wjf81ef <= tj8eafb;            ir7be3 <= qvabef4;            wwef8e7 <= fafbd2e;            ble39ca <= psf4b91;
         end      end
      generate         if ((twb8d6f==(plog2_points-2))&&(pdyn_points==1)) begin            assign jp4f44a = ui4cc50;            assign med12bd = qi3140a;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end         else if (twb8d6f==(plog2_points-1)) begin            assign jp4f44a = ui4cc50;            assign med12bd = qi3140a;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end         else if (pscale_reg==1) begin            assign jp4f44a = jp4acd7;            assign med12bd = swb35f0;            assign phbf55a = zz1cf94;            assign xwd56b8 = qi3e535;         end         else begin            assign jp4f44a = ui4cc50;            assign med12bd = qi3140a;            assign phbf55a = dmeb4a2;            assign xwd56b8 = bld2896;         end      endgenerate
      generate         if (pdyn_points==1) begin            if ((twb8d6f%2==0)&&(twb8d6f!=0)) begin                assign fn5ff31 = (hd940bd &(~qgeff2b)) | (vkb84a0 & qgeff2b) ;               assign eaff98f = (sj2f7f &(~qgeff2b)) | (rtc2502 & qgeff2b) ;               always @(negedge rstn or posedge clk) begin                  if (rstn==1'b0) begin                     dzc2d3f <= 'b0;                     wlb4ff7 <= 'b0;                  end                  else begin                                                               dzc2d3f <= qgeff2b ? {yx7f959[ks882e6-1],yx7f959[ks882e6-1:enc6b7b+1]} : hd2dec2;                     wlb4ff7 <= qgeff2b ? {yx7f959[enc6b7b-1],yx7f959[enc6b7b-1:1]} : xj7b0b4;
                  end               end               assign xy3fdeb = dzc2d3f;               assign shf7ad2 = wlb4ff7;
               always@(posedge clk or negedge rstn) begin	if(rstn==1'b0)	bl5f6cf<=0;	else	bl5f6cf <= aaacedc;               end               assign vifb67e = qgeff2b ? bl5f6cf : aaacedc;
            end            else if (twb8d6f%2==1) begin                assign fn5ff31 = hd940bd  ;               assign eaff98f = sj2f7f  ;               assign xy3fdeb = hd2dec2;               assign shf7ad2 = xj7b0b4;               assign vifb67e = aaacedc;            end            else begin               assign fn5ff31 = hd940bd  ;               assign eaff98f = sj2f7f  ;               assign xy3fdeb = hd2dec2;               assign shf7ad2 = xj7b0b4;               assign vifb67e=aaacedc;            end         end         else if ((twb8d6f%2==0)&&(twb8d6f!=0)) begin             assign fn5ff31 = hd940bd  ;            assign eaff98f = sj2f7f  ;            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  dzc2d3f <= 'b0;                  wlb4ff7 <= 'b0;               end               else begin                  dzc2d3f <= hd2dec2;                  wlb4ff7 <= xj7b0b4;               end            end            assign xy3fdeb = dzc2d3f;            assign shf7ad2 = wlb4ff7;
            assign vifb67e=aaacedc;         end         else begin            assign fn5ff31 = hd940bd  ;            assign eaff98f = sj2f7f  ;            assign xy3fdeb = hd2dec2;            assign shf7ad2 = xj7b0b4;
            assign vifb67e=aaacedc;         end      endgenerate
      generate         if ((pdyn_points==1)&&(twb8d6f<(plog2_points-2))) begin            assign gb4e6e8= lsbdfe5 ? {1'b0,uk2bfe6[hq35bdc-2:0]} : uk2bfe6[hq35bdc-1:0];         end         else if ((pdyn_points==0)&&(twb8d6f<(plog2_points-2))) begin            assign gb4e6e8= uk2bfe6;         end      endgenerate
         assign fnc8144     = pfdd15f;
         assign iccba1f = pffcacc[ks882e6-1:enc6b7b];      assign yxe87c3 = pffcacc[enc6b7b-1:0];
         assign wlbe0cb = wwe5667[vve6110-1:ptwid_widthr];      assign zm832e8 = wwe5667[ptwid_widthr-1:0];
         generate            if ((twb8d6f%2==0)&&(twb8d6f!=0))             osf5e4e_FFTC2048 # (               .hqadee3(hqadee3),               .pdin_widthr(enc6b7b),               .xj71cad(ptwid_widthr),               .plog2_points (plog2_points),               .xyadfc4(xyadfc4),               .phard_mac(phard_mac),               .device_family(med4d71)               )            ks15b47 (               .clk(clk),                         .rstn(rstn),                       .ph38443(iccba1f),                 .ri110f7(yxe87c3),                 .wlbe0cb(wlbe0cb),                   .zm832e8(zm832e8),                   .hbd80ed(hd2dec2),                 .ph3b7a(xj7b0b4)                  );         else if (twb8d6f%2==1) begin             assign gbf8740 = ic43e1d ? yxe87c3 : iccba1f;            assign cb1d024 = ic43e1d ? -iccba1f : yxe87c3;            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  nr4092d <= 'b0;                  sw24b7b <= 'b0;               end               else begin                  nr4092d <= gbf8740;                  sw24b7b <= cb1d024;               end            end             assign hd2dec2 = nr4092d;             assign xj7b0b4 = sw24b7b;
         end         else begin             assign hd2dec2 = iccba1f;             assign xj7b0b4 = yxe87c3;         end      endgenerate
         assign xl94d4c = dmeb4a2;      assign xy35331 = bld2896;      assign ui4cc50 = {xy3fdeb[enc6b7b-1],xy3fdeb};      assign qi3140a = {shf7ad2[enc6b7b-1],shf7ad2};
         assign vv50285 = xl94d4c + ui4cc50;      assign iea17e = xy35331 + qi3140a;      assign mt85f8e = xl94d4c - ui4cc50;      assign dz7e3ab = xy35331 - qi3140a;
               assign tj8eafb = {vv50285[ngb984-1],vv50285};      assign qvabef4 = {iea17e[ngb984-1],iea17e};      assign fafbd2e = {mt85f8e[ngb984-1],mt85f8e};      assign psf4b91 = {dz7e3ab[ngb984-1],dz7e3ab};
            generate         if((hqadee3==3)&&(twb8d6f%2==0)&&(twb8d6f!=0)) begin                   pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           shfd9c8 (            .clk               (clk),            .rstn              (rstn),            .din               (tj8eafb),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (ldfcc78),            .dout              (co2e45e)            );         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           ec824c5 (            .clk               (clk),            .rstn              (rstn),            .din               (qvabef4),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (the63c7),            .dout              (hd91781)            );         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           wl80422 (            .clk               (clk),            .rstn              (rstn),            .din               (fafbd2e),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (mg31e3e),            .dout              (cz5e07e)            );         pua7955_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           aab9f03 (            .clk               (clk),            .rstn              (rstn),            .din               (psf4b91),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (wl8f1f1),            .dout              (rv81fa0)            );
         end         else if (hqadee3==3) begin          yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           rg5843d (            .clk               (clk),            .rstn              (rstn),            .din               (tj8eafb),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (ldfcc78),            .dout              (co2e45e)            );         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           fc1b64c (            .clk               (clk),            .rstn              (rstn),            .din               (qvabef4),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (the63c7),            .dout              (hd91781)            );         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           ofc692e (            .clk               (clk),            .rstn              (rstn),            .din               (fafbd2e),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (mg31e3e),            .dout              (cz5e07e)            );         yzb4add_FFTC2048 #(            .twb8d6f       (twb8d6f),            .fc2aae9        (ngb984+1),            .epaba5f       (ngb984),            .fixed_scaling     (hqadee3),            .pdyn_points       (pdyn_points),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .plog2_points      (plog2_points),            .rounding_method   (rounding_method))           mta4b11 (            .clk               (clk),            .rstn              (rstn),            .din               (psf4b91),            .cz709f8             (vifb67e),            .qgeff2b            (qgeff2b),            .except            (wl8f1f1),            .dout              (rv81fa0)            );         end         else if((hqadee3==0)&&(twb8d6f%2==0)&&(twb8d6f!=0)) begin             assign co2e45e = {tj8eafb[ngb984-1],tj8eafb[ngb984-3+hqadee3:hqadee3],1'b0};            assign hd91781 = {qvabef4[ngb984-1],qvabef4[ngb984-3+hqadee3:hqadee3],1'b0};            assign cz5e07e = {fafbd2e[ngb984-1],fafbd2e[ngb984-3+hqadee3:hqadee3],1'b0};            assign rv81fa0 = {psf4b91[ngb984-1],psf4b91[ngb984-3+hqadee3:hqadee3],1'b0};
            assign ldfcc78= ^wjf81ef[ngb984-1:ngb984-2];            assign the63c7= ^ir7be3[ngb984-1:ngb984-2];            assign mg31e3e= ^wwef8e7[ngb984-1:ngb984-2];            assign wl8f1f1= ^ble39ca[ngb984-1:ngb984-2];         end         else if(hqadee3==0) begin             assign co2e45e = tj8eafb[ngb984-1+hqadee3:hqadee3];            assign hd91781 = qvabef4[ngb984-1+hqadee3:hqadee3];            assign cz5e07e = fafbd2e[ngb984-1+hqadee3:hqadee3];            assign rv81fa0 = psf4b91[ngb984-1+hqadee3:hqadee3];            assign ldfcc78= 1'b0;            assign the63c7= 1'b0;            assign mg31e3e= 1'b0;            assign wl8f1f1= 1'b0;         end      endgenerate
         assign jp7e838 = ipe8aff ? co2e45e : phbf55a;      assign dba0e32 = ipe8aff ? hd91781 : xwd56b8;      assign bn32d7d = ipe8aff ? cz5e07e : jp4f44a;      assign tjb5f73 = ipe8aff ? rv81fa0 : med12bd;      assign fp38cb5 = {jp7e838,dba0e32};
         assign kqff295 = {bn32d7d,tjb5f73};
      assign dmeb4a2 = go7dcff[wje829b-1:ngb984];      assign bld2896 = go7dcff[ngb984-1:0];
      generate      begin         if (twb8d6f==(plog2_points-1)) begin            assign go7dcff = neca54e;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-2))) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0)                  ks3b5bf <= 'b0;               else                  ks3b5bf <= neca54e;            end            assign go7dcff = lsbdfe5 ? neca54e : ks3b5bf;             end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==1)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  ks3b5bf  <= 'b0;                  mrd6fcb <= 'b0;                  phbf2ea <= 'b0;                  uicbabe <= 'b0;                  tu73fca  <= 'b0;               end               else begin                  ks3b5bf  <= neca54e;                  mrd6fcb <= ks3b5bf;                  phbf2ea <= mrd6fcb;                  uicbabe <= phbf2ea;                  tu73fca  <= lsbdfe5 ? kqff295 : ks3b5bf;               end            end            assign go7dcff = tu73fca;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==0)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0) begin                  ks3b5bf  <= 'b0;                  mrd6fcb <= 'b0;                  phbf2ea <= 'b0;                  uicbabe <= 'b0;                  tu73fca  <= 'b0;               end               else begin                  ks3b5bf  <= neca54e;                  mrd6fcb <= ks3b5bf;                  phbf2ea <= mrd6fcb;                  uicbabe <= phbf2ea;                  tu73fca  <= lsbdfe5 ? neca54e : mrd6fcb;               end            end            assign go7dcff = tu73fca;         end         else if ((pdyn_points==0)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==1)) begin            assign go7dcff = neca54e;         end         else if ((pdyn_points==0)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==0)) begin            always @(negedge rstn or posedge clk) begin               if (rstn==1'b0)                  ks3b5bf <= 'b0;               else                  ks3b5bf <= neca54e;            end            assign go7dcff = ks3b5bf;         end         else begin            me5334a_FFTC2048 #(               .ba99a50(wje829b),               .ho69416(hq35bdc),               .gq1a9ae(gq1a9ae),               .med4d71(med4d71)               )           qv9fe30 (               .clk(clk),                        .rstn(rstn),                      .pfdd15f(pfdd15f),                    .uk2bfe6(gb4e6e8),                 .neca54e(neca54e),                  .tj9ba2b(tj9ba2b),                    .go7dcff(go7dcff)                 );         end      end      endgenerate
         ea78733_FFTC2048 #(         .pdyn_points  (pdyn_points),         .plog2_points (plog2_points),         .twb8d6f  (twb8d6f),         .yz26d41  (hq35bdc),         .xlb506c  (xj7b8d4),         .ip41b33 (bn2219e),         .pscale_reg   (pscale_reg),         .fc3fcb5(fc3fcb5),         .gq1a9ae(gq1a9ae)         )      rg5282c (            .clk(clk),                     .rstn(rstn),                   .mt12817    (mt12817),             .qi5137(qi5137),                     .lsbdfe5(lsbdfe5),            .hd940bd(fn5ff31),               .tja05ef(tja05ef),               .sj2f7f(eaff98f),               .qv17bfc(qv17bfc),               .os67205(os67205),            .ipe8aff(ipe8aff),                   .ic43e1d(ic43e1d),               .pfdd15f(pfdd15f),                 .uk2bfe6(uk2bfe6),                 .tj9ba2b(tj9ba2b),                 .bn289b8(bn289b8)                  );
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            en44dc6 <= 'b0;            neca54e <= 'b0;         end         else begin            en44dc6 <= fp38cb5;            neca54e <= kqff295;         end      end
      generate         if (twb8d6f==(plog2_points-1)) begin            assign vif1a71 = fn5ff31;         end         else  begin            assign vif1a71 = encce40;         end      endgenerate
      generate         if ((pdyn_points==1)&&(vv7105c==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  an39028 <= 1'b1;               end               else begin                  if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                                       an39028 <= ~an39028;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  zxc7c69 <= 1'b0;               end               else begin                                                      if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                     zxc7c69 <= 1'b0;                                    else if (ou8d38b)                     zxc7c69 <= zxc7c69 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                                                      if (((vif1a71)||(cm599c8))&&(an39028==ou2b339))                     vv40a26 <= 1'b0;                  else if (an39028==ou2b339)                     vv40a26 <= zxc7c69;               end            end
         end         else if ((pdyn_points==0)&&(vv7105c==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  an39028 <= 1'b1;               end               else begin                  if (vif1a71)                     an39028 <= ~an39028;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  zxc7c69 <= 1'b0;               end               else begin                  if (vif1a71)                     zxc7c69 <= 1'b0;                                    else if (ou8d38b)                     zxc7c69 <= zxc7c69 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                  if (vif1a71)                     vv40a26 <= 1'b0;                  else if (an39028==ou2b339)                     vv40a26 <= zxc7c69;               end            end
         end         else begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  vv40a26 <= 1'b0;               end               else begin                  if (vif1a71)                     vv40a26 <= 1'b0;                                    else if (ou8d38b)                     vv40a26 <= vv40a26 | ldfcc78 | the63c7 | mg31e3e | wl8f1f1;               end            end        end     endgenerate
   endmodule                                                                                                   
`timescale 1 ns / 100 ps
module me5334a_FFTC2048 (
            clk,       
            rstn,      
            pfdd15f,     
            uk2bfe6,     
            neca54e,    
            tj9ba2b,     
            go7dcff    
            );
parameter ba99a50      = 16;
parameter ho69416      = 16;
parameter gq1a9ae     = 1;
parameter med4d71 = "ECP";
localparam kqde610   = 1<<ho69416;
input                      clk;
input                      rstn;
input                      pfdd15f;
input  [ho69416-1:0]     uk2bfe6;
input  [ba99a50-1:0]     neca54e;
input  [ho69416-1:0]     tj9ba2b;
output [ba99a50-1:0]     go7dcff;
reg    [ba99a50-1:0]     uv5be0e;
wire   [ba99a50-1:0]     alf83aa;
wire                       cmc1d54;
wire                       vkeaa1;
reg    [ba99a50-1:0]     phaa854;
                                          assign cmc1d54 = 1'b1;      assign vkeaa1 = 1'b1;
      generate
      if (gq1a9ae==0) begin         pmi_distributed_dpram  #(            .pmi_addr_depth         (kqde610),            .pmi_addr_width         (ho69416),            .pmi_data_width         (ba99a50),            .pmi_regmode            ("reg"),            .pmi_init_file          ("none"),            .pmi_init_file_format   ("binary"),            .pmi_family             (med4d71),            .module_type            ("pmi_distributed_dpram")            )            ea688fd (               .WrAddress   (uk2bfe6),               .Data        (neca54e),               .WrClock     (clk),               .WE          (pfdd15f),               .WrClockEn   (vkeaa1),               .RdAddress   (tj9ba2b),               .RdClock     (clk),               .RdClockEn   (cmc1d54),               .Reset       (~rstn),               .Q           (alf83aa)               );
         assign go7dcff = alf83aa;
      end      else begin         pmi_ram_dp #(            .pmi_wr_addr_depth         (kqde610),            .pmi_wr_addr_width         (ho69416),            .pmi_wr_data_width         (ba99a50),            .pmi_rd_addr_depth         (kqde610),            .pmi_rd_addr_width         (ho69416),            .pmi_rd_data_width         (ba99a50),            .pmi_gsr                   ("disable"),            .pmi_resetmode             ("sync"),            .pmi_init_file             ("none"),            .pmi_init_file_format      ("binary"),            .pmi_regmode               ("reg"),            .pmi_family                (med4d71),            .module_type               ("pmi_ram_dp")            )         ui536e7 (               .WrAddress   (uk2bfe6),               .RdAddress   (tj9ba2b),               .Data        (neca54e),               .RdClock     (clk),               .WrClock     (clk),               .RdClockEn   (cmc1d54),               .WrClockEn   (vkeaa1),               .WE          (pfdd15f),               .Reset       (1'b0),               .Q           (alf83aa)               );
            always @(posedge clk or negedge rstn) begin            if(rstn==1'b0)               uv5be0e <= 'b0;            else               uv5be0e <= alf83aa;         end
         assign go7dcff = uv5be0e;      end
      endgenerate
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module aabcb24_FFTC2048 (
              clk,               
              rstn,              
              fft_mode,          
              ec24226,            
              dire,              
              diim,              
              dore,              
              doim               
              ) ;
parameter fc2aae9   = 16;
parameter ls89b60   = 1;
input                      clk;
input                      rstn;
input                      fft_mode ;
input                      ec24226;
input [fc2aae9-1:0]     dire;
input [fc2aae9-1:0]     diim;
output [fc2aae9-1:0]    dore;
output [fc2aae9-1:0]    doim;
reg [fc2aae9-1:0]       dore;
reg [fc2aae9-1:0]       doim;
                        generate          if (ls89b60==1) begin                            always @(posedge clk or negedge rstn)              begin                 if(!rstn)                    doim <= {fc2aae9{1'b0}};                 else begin                    if(ec24226==1'b1)	doim <= fft_mode ? (1'b1 + (~diim)) : diim;                    else	doim <= 'b0;                 end              end
                            always @(posedge clk or negedge rstn)              begin                 if(!rstn) dore <= {fc2aae9{1'b0}};                 else begin                    if(ec24226==1'b1)	dore <= dire; else	dore <= 'b0;                 end              end          end          else begin                              always @(posedge clk or negedge rstn)              begin                 if(!rstn)                    doim <= {fc2aae9{1'b0}};                 else                    doim <= fft_mode ? (1'b1 + (~diim)) : diim;              end
                            always @(posedge clk or negedge rstn)              begin                 if(!rstn)                    dore <= {fc2aae9{1'b0}};                 else dore <= dire;              end          end      endgenerate   endmodule                                                                                             
`timescale 1 ns / 100 ps
module ea78733_FFTC2048 (
            clk,       
            rstn,      
            mt12817,     
            lsbdfe5, 
            hd940bd,    
            tja05ef,    
            sj2f7f,    
            qv17bfc,    
            os67205,  
            qi5137,       
            ipe8aff,      
            ic43e1d,    
            pfdd15f,     
            uk2bfe6,     
            tj9ba2b,     
            bn289b8      
            ) ;
parameter pdyn_points  = 0;
parameter plog2_points = 4;
parameter twb8d6f  = 0;
parameter yz26d41  = 4;
parameter xlb506c  = 4;
parameter ip41b33 = 1;
parameter gq1a9ae   = 1;
parameter pscale_reg   = 0;
parameter fc3fcb5 = 3;
localparam rib864c         = (1<<plog2_points)-1;
localparam jr19315      = (1<<yz26d41)-4;
localparam ay4c57d      = (1<<yz26d41)-3;
localparam aa15f41         = (1<<yz26d41)-2;
localparam ic7d047          = (gq1a9ae==0) ? ay4c57d : jr19315;
localparam by47165           = (twb8d6f%2==0)?1:0;
localparam xwc595f          = (twb8d6f%2==1)?1:0;
localparam ip657dc          = (1<<yz26d41);
localparam xj5f729          = (twb8d6f%2==0)?(ip657dc+1):(ip657dc+fc3fcb5);
localparam al4e50c          = ip657dc-6;
localparam nt94328         = plog2_points+1-twb8d6f;
localparam sh651e7        = plog2_points-1-twb8d6f;
localparam qv3cf72         = twb8d6f-2;
localparam tj3dcad     = nt94328  -1;
localparam su72b7a    = sh651e7 -1;
localparam riade84     = qv3cf72  +1;
localparam mr7a114          = (3*ip657dc)-3;
localparam db8452a            = (4*ip657dc)-3;
localparam do14ab7     = (pscale_reg==1) ? (1<<plog2_points)-7 : (1<<plog2_points)-6;
localparam vkb75d9       = (1<<(yz26d41-1));
localparam ldd765e     = ic7d047 - vkb75d9;
localparam iccbdad    = aa15f41 - vkb75d9;
localparam fpb5a2e     = xj5f729 - vkb75d9;
localparam dz45dd8 = xj5f729 - vkb75d9 - 2;
localparam mtbb1c9      = (1<<(yz26d41-1));
localparam xjc726e     = (3*mtbb1c9)-3;
localparam qtc9bbc       = (4*mtbb1c9)-3;
localparam pf6ef2b     = mtbb1c9-6;
input                      clk;
input                      rstn;
input  [plog2_points-1:0]  mt12817;
input                      hd940bd;
input                      sj2f7f;
input                      lsbdfe5;
output                     tja05ef;
output                     qv17bfc;
output                     os67205;
output                     qi5137;
output                     ipe8aff;
output                     ic43e1d;
output                     pfdd15f;
output  [plog2_points-1:0] uk2bfe6;
output  [yz26d41-1:0]  tj9ba2b;
output  [xlb506c-1:0]  bn289b8;
reg     [plog2_points-1:0] hbe306d ;
reg                        wl1836e ;
wire                       qi5137 ;
reg     [yz26d41-1:0]  ui6dd4d ;
reg                        bl6ea68;
wire                       ip75347;
wire                       ksa9a3c;
reg                        xw4d1e0;
reg                        go68f02;
reg     [plog2_points-1:0] ir3c082;
reg     [plog2_points-1:0] bn289b8;
wire    [nt94328+1:0]  ou82869;
wire    [nt94328+1:0]  ira1a43;
reg                        epd21c ;
wire                       lq690e4 ;
reg     [plog2_points-1:0] yk4391a;
reg     [plog2_points-1:0] nee4686;
reg     [plog2_points-1:0] ks1a19c;
wire                       hd940bd;
reg                        zm86702;
reg                        yz33813;
wire                       tja05ef;
wire                       kqe04e3;
wire                       yz2719;
wire                       rv138cd;
reg                        tw9c66f;
reg                        pfe337b;
wire                       sj2f7f;
reg                        jpcdef6;
reg                        en6f7b7;
reg                        dz7bdbc;
reg                        aydede6;
wire                       ipe8aff;
reg                        os67205;
reg                        ksbcc72;
reg                        lde6391;
reg                        aa31c8e;
reg                        ic43e1d;
reg                        ww7238f;
reg                        zz91c79;
wire  [plog2_points-1:0]   jp71e77;
wire  [plog2_points-1:0]   tu79dfd;
wire  [plog2_points-2:0]   ui77f58;
wire  [plog2_points-2:0]   shfd606;
wire  [yz26d41-1:0]    by581a2;
wire  [plog2_points-1:0]   zz689b;
wire  [plog2_points-1:0]   nga26f0;
wire  [yz26d41-1:0]    hd9bc16;
wire  [plog2_points+1:0]   qgf05b8;
wire  [plog2_points+1:0]   xl16e00;
wire  [plog2_points-2:0]   twb803b;
wire                       zkc01da;
wire                       swed2;
wire  [yz26d41+1:0]    ie3b48d;
reg                        tuda469;
                                    
            
                                                                                       generate      begin         if ((pdyn_points==1)&&(twb8d6f<(plog2_points-1))&&(twb8d6f%2==0)&&(twb8d6f!=0)) begin             assign ou82869={1'b0,ir3c082[sh651e7:0],1'b0}+{2'b0,ir3c082[sh651e7:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ks1a19c <= 'b0;               end               else begin                  case(ir3c082[nt94328:nt94328-1])                     2'b00: ks1a19c <='b0;                      2'b01: ks1a19c <=({ir3c082[sh651e7:0],1'b0})<<qv3cf72;                      2'b10: ks1a19c <=(ir3c082[sh651e7:0])<<qv3cf72;                      2'b11: ks1a19c <=(ou82869)<<qv3cf72;                   endcase               end            end            assign ira1a43={1'b0,ir3c082[su72b7a:0],1'b0}+{2'b0,ir3c082[su72b7a:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  nee4686 <= 'b0;               end               else begin                  case(ir3c082[tj3dcad:tj3dcad-1])                     2'b00: nee4686 <='b0;                      2'b01: nee4686 <=({ir3c082[su72b7a:0],1'b0})<<riade84;                      2'b10: nee4686 <=(ir3c082[su72b7a:0])<<riade84;                      2'b11: nee4686 <=(ira1a43)<<riade84;                   endcase               end            end            always @(*) begin               if (lsbdfe5)                  bn289b8 = nee4686;               else                  bn289b8 = ks1a19c;            end         end         else if ((pdyn_points==1)&&(twb8d6f%2==0)&&(twb8d6f==(plog2_points-1))) begin            assign ou82869={1'b0,ir3c082[sh651e7:0],1'b0}+{2'b0,ir3c082[sh651e7:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  bn289b8 <= 'b0;               end               else begin                  case(ir3c082[nt94328:nt94328-1])                     2'b00: bn289b8 <='b0;                      2'b01: bn289b8 <=({ir3c082[sh651e7:0],1'b0})<<qv3cf72;                      2'b10: bn289b8 <=(ir3c082[sh651e7:0])<<qv3cf72;                      2'b11: bn289b8 <=(ou82869)<<qv3cf72;                   endcase               end            end         end         else if ((pdyn_points==0)&&(twb8d6f%2==0)&&(twb8d6f!=0)) begin            assign ou82869={1'b0,ir3c082[sh651e7:0],1'b0}+{2'b0,ir3c082[sh651e7:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  bn289b8 <= 'b0;               end               else begin                  case(ir3c082[nt94328:nt94328-1])                     2'b00: bn289b8 <='b0;                      2'b01: bn289b8 <=({ir3c082[sh651e7:0],1'b0})<<qv3cf72;                      2'b10: bn289b8 <=(ir3c082[sh651e7:0])<<qv3cf72;                      2'b11: bn289b8 <=(ou82869)<<qv3cf72;                   endcase               end            end         end      end      endgenerate
         generate      begin         if (pdyn_points==1) begin            assign jp71e77     = mt12817;            assign ui77f58      = lsbdfe5 ? ldd765e  :ic7d047 ;            assign shfd606     = lsbdfe5 ? iccbdad :aa15f41 ;            assign zz689b      = lsbdfe5 ? fpb5a2e :xj5f729 ;            assign nga26f0  = lsbdfe5 ? dz45dd8: xj5f729;            assign qgf05b8      = lsbdfe5 ? xjc726e :mr7a114 ;            assign xl16e00        = lsbdfe5 ? qtc9bbc :db8452a ;            assign twb803b      = lsbdfe5 ? pf6ef2b :al4e50c ;            assign zkc01da = hd940bd;            assign swed2 = sj2f7f;         end         else begin            assign jp71e77     = rib864c;            assign ui77f58      = ic7d047;            assign shfd606     = aa15f41;            assign zz689b      = xj5f729;            assign nga26f0  = xj5f729;            assign qgf05b8      = mr7a114 ;            assign xl16e00        = db8452a ;            assign twb803b      = al4e50c ;            assign zkc01da = 1'b0;            assign swed2 = 1'b0;         end      end      endgenerate
      generate      begin         if ((pdyn_points==1)&&(pscale_reg==0)) begin            assign tu79dfd = mt12817 - 5;            assign rv138cd    = lde6391;         end         else if ((pdyn_points==1)&&(pscale_reg==1)) begin            assign tu79dfd = mt12817 - 6;            assign rv138cd    = aa31c8e;         end         else begin            assign tu79dfd = do14ab7 ;            assign rv138cd    = lde6391;         end      end      endgenerate
         generate      begin         if ((pdyn_points==1)&&(yz26d41>1)) begin            assign by581a2      = lsbdfe5 ? uk2bfe6[yz26d41-2:0] :uk2bfe6[yz26d41-1:0] ;            assign hd9bc16  = lsbdfe5 ? {1'b0,ui6dd4d[yz26d41-2:0]} :ui6dd4d ;         end         else if ((pdyn_points==1)&&(yz26d41==1)) begin            assign by581a2      = uk2bfe6[yz26d41-1:0] ;            assign hd9bc16  = lsbdfe5 ? {1'b0,ui6dd4d[yz26d41-1:0]} :ui6dd4d ;         end         else if (pdyn_points==0) begin            assign hd9bc16  = ui6dd4d ;         end      end      endgenerate
         generate      begin         if ((gq1a9ae==0)&&(pscale_reg==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  tuda469 <= 1'b0;               end               else begin                  tuda469 <= ((hbe306d==(ui77f58-1))&&(wl1836e)) ? 1'b1 : 1'b0;               end            end         end         else if ((gq1a9ae>0)&&(pscale_reg==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  tuda469 <= 1'b0;               end               else begin                  tuda469 <= ((hbe306d==(ui77f58-2))&&(wl1836e)) ? 1'b1 : 1'b0;               end            end         end         else if ((gq1a9ae==0)&&(pscale_reg==1)&&(twb8d6f==(plog2_points-4))&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  tuda469 <= 1'b0;               end               else begin                  if (lsbdfe5)                     tuda469 <= hd940bd;                  else                     tuda469 <= ((hbe306d==(ui77f58-2))&&(wl1836e)) ? 1'b1 : 1'b0;               end            end         end         else if ((gq1a9ae==0)&&(pscale_reg==1)&&(twb8d6f==(plog2_points-3))) begin            always @(*) begin                  tuda469 = zm86702;            end         end         else if ((gq1a9ae==0)&&(pscale_reg==1)&&(twb8d6f!=(plog2_points-3))) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  tuda469 <= 1'b0;               end               else begin                  tuda469 <= ((hbe306d==(ui77f58-2))&&(wl1836e)) ? 1'b1 : 1'b0;               end            end         end         else if ((gq1a9ae>0)&&(pscale_reg==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  tuda469 <= 1'b0;               end               else begin                  tuda469 <= ((hbe306d==(ui77f58-3))&&(wl1836e)) ? 1'b1 : 1'b0;               end            end         end      end      endgenerate
                  always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            hbe306d <= 'b0;         else if (zkc01da==1'b1)            hbe306d <= 'b0;         else if (wl1836e==1'b1)            hbe306d <= hbe306d+1;      end
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            wl1836e <= 1'b0;         else if (hd940bd==1'b1)            wl1836e <= 1'b1;         else if (qi5137==1'b1)            wl1836e <= 1'b0;      end
         assign qi5137 = (hbe306d==jp71e77)? 1'b1 : 1'b0;
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            ui6dd4d <= 'b0;         else if (ksa9a3c==1'b1)            ui6dd4d <= 'b0;         else if (bl6ea68)            ui6dd4d <= ui6dd4d+1;      end
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            bl6ea68 <= 1'b0;         else if (ksa9a3c==1'b1)            bl6ea68 <= 1'b1;         else if (ip75347==1'b1)            bl6ea68 <= 1'b0;      end
         assign ip75347 = (hd9bc16==jp71e77)? 1'b1 : 1'b0;
         assign ksa9a3c = tuda469;
            generate         if ((twb8d6f%2==0)&&(twb8d6f!=0)) begin                         always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  epd21c <= 1'b0;               else if (sj2f7f==1'b1)                  epd21c <= 1'b1;               else if (lq690e4==1'b1)                  epd21c <= 1'b0;            end                        assign lq690e4 = (ir3c082==jp71e77)? 1'b1 : 1'b0;            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ir3c082 <= 'b0;               else if (swed2==1'b1)                  ir3c082 <= 'b0;               else if (epd21c==1'b1)                  ir3c082 <= ir3c082+1;            end         end      endgenerate
      always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            zm86702  <= 1'b0;            yz33813 <= 1'b0;            aydede6   <= 1'b0;            tw9c66f   <= 1'b0;            pfe337b   <= 1'b0;         end         else begin            zm86702  <= hd940bd;            yz33813 <= zm86702;            aydede6   <= dz7bdbc;            tw9c66f   <= kqe04e3;            pfe337b   <= yz2719;         end      end            always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ksbcc72  <= 1'b0;            lde6391 <= 1'b0;            aa31c8e <= 1'b0;         end         else  begin            ksbcc72  <= os67205;            lde6391 <= ksbcc72;            aa31c8e <= lde6391;         end      end            always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            ww7238f <= 1'b0;         else if (hd940bd)            ww7238f <= 1'b1;         else if (rv138cd)            ww7238f <= 1'b0;      end
         generate      begin         if ((pdyn_points==1)&&(twb8d6f==(plog2_points-1))) begin                           assign kqe04e3 = zm86702;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-2))&&(twb8d6f%2==1)) begin               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= lsbdfe5 ? hd940bd: ((hbe306d==(zz689b)) ? 1'b1 : 1'b0);            end            assign kqe04e3 = lsbdfe5 ? zm86702: ((hbe306d==(zz689b+1)) ? 1'b1 : 1'b0);                     end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-2))) begin               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= lsbdfe5 ? hd940bd: ((hbe306d==(zz689b-1)) ? 1'b1 : 1'b0);            end            assign kqe04e3 = lsbdfe5 ? zm86702: ((hbe306d==(zz689b)) ? 1'b1 : 1'b0);                     end         else if ((pdyn_points==1)&&(twb8d6f<(plog2_points-2))&&(twb8d6f%2==1)) begin               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= (hbe306d==zz689b) ? 1'b1 : 1'b0;            end            assign kqe04e3 = (hbe306d==(zz689b+1)) ? 1'b1 : 1'b0;         end         else if ((pdyn_points==1)&&(twb8d6f<(plog2_points-2))) begin               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= (hbe306d==(zz689b-1)) ? 1'b1 : 1'b0;            end            assign kqe04e3 = (hbe306d==zz689b) ? 1'b1 : 1'b0;         end         else if ((pdyn_points==0)&&(twb8d6f==(plog2_points-1))) begin               assign kqe04e3 = zm86702;         end         else if ((pdyn_points==0)&&(twb8d6f<(plog2_points-1))&&(twb8d6f%2==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= (hbe306d==xj5f729) ? 1'b1 : 1'b0;            end            assign kqe04e3 = zz91c79;         end         else if ((pdyn_points==0)&&(twb8d6f<(plog2_points-1))) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  zz91c79 <= 1'b0;               else                  zz91c79 <= (hbe306d==(xj5f729-1)) ? 1'b1 : 1'b0;            end            assign kqe04e3 = zz91c79;         end      end      endgenerate         generate         if((pdyn_points==1)&&(plog2_points%2==1)&&(xwc595f==1)&&(twb8d6f==(plog2_points-4))&&(pscale_reg==1))  begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  jpcdef6  <= 1'b0;               end               else begin                  jpcdef6  <= sj2f7f;               end            end            assign yz2719 = lsbdfe5 ? jpcdef6 : ((hbe306d==twb803b) ? 1'b1 : 1'b0);         end         else if((pdyn_points==1)&&(plog2_points%2==1)&&(xwc595f==1)&&(twb8d6f==(plog2_points-4))&&(pscale_reg==0))            assign yz2719 = lsbdfe5 ? sj2f7f : ((hbe306d==twb803b) ? 1'b1 : 1'b0);         else if((xwc595f==1)&&(twb8d6f<(plog2_points-3)))             assign yz2719 = (hbe306d==twb803b) ? 1'b1 : 1'b0;         else if((pdyn_points==1)&&(plog2_points%2==1)&&(by47165==1)&&(twb8d6f==(plog2_points-5)))            assign yz2719 = (hbe306d==(nga26f0+1)) ? 1'b1 : 1'b0;         else if((xwc595f==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==0))             assign yz2719 = sj2f7f;         else if((xwc595f==1)&&(twb8d6f==(plog2_points-3))&&(pscale_reg==1)) begin             always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  jpcdef6  <= 1'b0;               end               else begin                  jpcdef6  <= sj2f7f;               end            end            assign yz2719 = jpcdef6;         end         else if((xwc595f==1)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==0))             assign yz2719 = sj2f7f;         else if((xwc595f==1)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==1)&&(pdyn_points==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  jpcdef6  <= 1'b0;                  en6f7b7 <= 1'b0;               end               else begin                  jpcdef6   <= sj2f7f;                  en6f7b7  <= jpcdef6;               end            end            assign yz2719 = en6f7b7;         end         else if((xwc595f==1)&&(twb8d6f==(plog2_points-2))&&(pscale_reg==1)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  jpcdef6  <= 1'b0;                  en6f7b7 <= 1'b0;               end               else begin                  jpcdef6   <= sj2f7f;                  en6f7b7  <= jpcdef6;               end            end            assign yz2719 = jpcdef6;         end         else if((by47165==1)&&(twb8d6f==(plog2_points-4)))             assign yz2719 = (hbe306d==(nga26f0-1)) ? 1'b1 : 1'b0;         else if((by47165==1)&&(twb8d6f==(plog2_points-3))) begin             always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  xw4d1e0  <= 1'b0;                  go68f02 <= 1'b0;               end               else begin                  xw4d1e0  <= ksa9a3c;                  go68f02 <= xw4d1e0;               end            end            assign yz2719 = xw4d1e0;         end         else            assign yz2719 = 1'b0;      endgenerate
               generate                                                               if ((pdyn_points==1)&&(pscale_reg==1)&&(twb8d6f!=(plog2_points-3))&&(twb8d6f!=(plog2_points-2))&&(twb8d6f!=(plog2_points-1))) begin            assign ipe8aff = dz7bdbc;            assign tja05ef = tw9c66f;            assign qv17bfc = yz2719;         end         else if ((pdyn_points==1)&&(pscale_reg==1)&&((twb8d6f==(plog2_points-3))||(twb8d6f==(plog2_points-2))||(twb8d6f!=(plog2_points-1)))) begin            assign ipe8aff = dz7bdbc;            assign tja05ef = kqe04e3;            assign qv17bfc = yz2719;         end         else if ((pscale_reg==1)&&(twb8d6f!=(plog2_points-2))&&(twb8d6f!=(plog2_points-1))) begin            assign ipe8aff = dz7bdbc;            assign tja05ef = tw9c66f;            assign qv17bfc = yz2719;         end         else if ((pscale_reg==1)&&((twb8d6f==(plog2_points-2))||(twb8d6f!=(plog2_points-1)))) begin            assign ipe8aff = dz7bdbc;            assign tja05ef = kqe04e3;            assign qv17bfc = yz2719;         end         else if ((pdyn_points==1)&&(twb8d6f==(plog2_points-1))) begin            assign ipe8aff = lsbdfe5 ? 1'b0 : dz7bdbc;            assign tja05ef = kqe04e3;            assign qv17bfc = yz2719;         end         else begin            assign ipe8aff = dz7bdbc;            assign tja05ef = kqe04e3;            assign qv17bfc = yz2719;         end      endgenerate
      generate      begin         if ((pdyn_points==1)&&(yz26d41>1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  dz7bdbc <= 1'b0;               else if (hd940bd==1'b1)                  dz7bdbc <= 1'b0;               else if ((by581a2[yz26d41-1:0]==shfd606)&&(wl1836e))                  dz7bdbc <= ~dz7bdbc;            end         end         else if ((pdyn_points==1)&&(yz26d41==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  dz7bdbc <= 1'b0;               else if (lsbdfe5==1'b1) begin                  if (hd940bd)                     dz7bdbc <= ~dz7bdbc;                  else if (qi5137==1'b1)                     dz7bdbc <= 1'b0;                  else if (wl1836e)                     dz7bdbc <= ~dz7bdbc;               end               else if (hd940bd==1'b1)                  dz7bdbc <= 1'b0;               else if ((by581a2[0:0]==shfd606)&&(wl1836e))                  dz7bdbc <= ~dz7bdbc;            end         end         else if ((pdyn_points==0)&&(yz26d41>0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  dz7bdbc <= 1'b0;               else if (hd940bd==1'b1)                  dz7bdbc <= 1'b0;               else if ((uk2bfe6[yz26d41-1:0]==aa15f41)&&(wl1836e))                  dz7bdbc <= ~dz7bdbc;            end         end         else begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  dz7bdbc <= 1'b0;               else if (hd940bd)                  dz7bdbc <= ~dz7bdbc;               else if (qi5137==1'b1)                  dz7bdbc <= 1'b0;               else if (wl1836e)                  dz7bdbc <= ~dz7bdbc;            end         end      end      endgenerate
         generate      begin         if ((pdyn_points==1)&&((xwc595f==1)&&(twb8d6f<(plog2_points-1)))&&(pscale_reg==0)) begin            assign ie3b48d = {(uk2bfe6[yz26d41+1]&(~lsbdfe5)),uk2bfe6[yz26d41:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if (ww7238f) begin                  if (ie3b48d==qgf05b8)                     ic43e1d <= 1'b1;                  else if (ie3b48d==xl16e00)                     ic43e1d <= 1'b0;               end            end         end         else if ((pdyn_points==1)&&((xwc595f==1)&&(twb8d6f<(plog2_points-2)))&&(pscale_reg==1)) begin            assign ie3b48d = {(uk2bfe6[yz26d41+1]&(~lsbdfe5)),uk2bfe6[yz26d41:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if (ww7238f) begin                  if (ie3b48d==(qgf05b8-1))                     ic43e1d <= 1'b1;                  else if (ie3b48d==(xl16e00-1))                     ic43e1d <= 1'b0;               end            end         end         else if ((pdyn_points==1)&&((xwc595f==1)&&(twb8d6f==(plog2_points-2)))&&(pscale_reg==1)) begin            assign ie3b48d = {(uk2bfe6[yz26d41+1]&(~lsbdfe5)),uk2bfe6[yz26d41:0]};            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if (ww7238f) begin                  if (ie3b48d==qgf05b8)                     ic43e1d <= 1'b1;                  else if (ie3b48d==xl16e00)                     ic43e1d <= 1'b0;               end            end         end         else if ((pdyn_points==0)&&((xwc595f==1)&&(twb8d6f<(plog2_points-1)))&&(pscale_reg==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if (uk2bfe6[yz26d41+1:0]==mr7a114)                  ic43e1d <= 1'b1;               else if (uk2bfe6[yz26d41+1:0]==db8452a)                  ic43e1d <= 1'b0;            end         end         else if ((pdyn_points==0)&&((xwc595f==1)&&(twb8d6f<(plog2_points-1)))&&(pscale_reg==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if (uk2bfe6[yz26d41+1:0]==(mr7a114-1))                  ic43e1d <= 1'b1;               else if (uk2bfe6[yz26d41+1:0]==(db8452a-1))                  ic43e1d <= 1'b0;            end         end         else if((xwc595f==1)&&(twb8d6f==(plog2_points-1)))             always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  ic43e1d <= 1'b0;               else if ((uk2bfe6[1:0]==2'b0)&&(wl1836e==1'b1))                  ic43e1d <= 1'b1;               else                  ic43e1d <= 1'b0;            end      end      endgenerate
         assign pfdd15f = wl1836e;      assign uk2bfe6 = hbe306d;      generate         if(twb8d6f==(plog2_points-2))             assign tj9ba2b = uk2bfe6;         else            assign tj9ba2b = hd9bc16[yz26d41-1:0];      endgenerate
         
   always @(posedge clk or negedge rstn)   begin      if(!rstn)         os67205 <= 1'b0;      else         os67205 <= (hbe306d==tu79dfd)? 1'b1 : 1'b0;   end
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module wwdbe0f_FFTC2048 (
                clk,       
                rstn,      
                mec1e54,   
                ibstart,   
                os67205,  
                qi5137,       
                of54252,   
                wla1295,
                rv94ad, 
                cm599c8,  
                jc52b77, 
                ir95bbb, 
                ibend,     
                rfib       
                );
parameter bit_reverse   = 0;
parameter pdyn_points   = 0;
input                        clk;
input                        rstn;
input                        mec1e54;
input                        ibstart;
input                        os67205;
input                        qi5137;
input                        of54252;
input                        jc52b77;
input                        rv94ad;
input                        cm599c8;
input                        wla1295;
output                       ir95bbb;
output                       ibend;
output                       rfib;
reg                          ibend;
reg                          rfib;
reg                          tu529c6;
reg                          lf94e33;
reg                          twa719e;
reg                          ph38cf2;
reg                          yxc6797;
reg                          qv33cbd;
reg                          zz9e5ec;
reg                          gbf2f66;
reg                          uk97b34;
reg                          ribd9a1;
wire                         pfecd0b;
reg                          lq6685e;
reg	ec342f3;
reg [2:0]	gda1798;
reg [2:0]	ribcc5;
wire	mr5e62a;
            
                     generate         if ((bit_reverse==0) || ((bit_reverse==1)&&(pdyn_points==0))) begin              always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  qv33cbd  <= 1'b0;               end               else begin                  if (rv94ad)                     qv33cbd <= yxc6797;               end            end         end         else if (pdyn_points==1)  begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  qv33cbd  <= 1'b0;               end               else begin                  if (cm599c8)                     qv33cbd <= yxc6797;               end            end         end      endgenerate
      always@(posedge clk or negedge rstn) begin         if(rstn==1'b0)	ec342f3 <=1'b0;         else if(ibstart)	ec342f3 <= 1'b1;      end
      generate         if (bit_reverse==0) begin              assign pfecd0b      = ec342f3 ? of54252 : 1'b0;            assign ir95bbb = zz9e5ec;         end         else begin            assign ir95bbb = qv33cbd;            assign pfecd0b      = ec342f3 ? qi5137 : 1'b0;         end      endgenerate
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ibend    <= 1'b0;            tu529c6  <= 1'b1;            lf94e33  <= 1'b1;            twa719e  <= 1'b0;            ph38cf2  <= 1'b0;            yxc6797  <= 1'b0;            zz9e5ec  <= 1'b0;            ribd9a1     <= 1'b0;         end         else begin            ribd9a1     <= ibstart;            if (os67205)               ibend <= 1'b1;            else               ibend <= 1'b0;            tu529c6  <= rfib;            lf94e33  <= tu529c6;            if (ph38cf2)               yxc6797 <= jc52b77;            if (cm599c8)               zz9e5ec <= qv33cbd;            twa719e  <= os67205;            ph38cf2  <= twa719e;         end      end
         generate      begin         if (pdyn_points==0) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  rfib     <= 1'b1;               end               else begin                  if (os67205)                     rfib <= 1'b1;                  else if (ibstart&&lf94e33)                     rfib <= 1'b0;               end            end         end         else  begin                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            always @(posedge clk or negedge rstn) begin	if(rstn==1'b0) begin	gda1798<=0;	end	else begin	if(mec1e54)	gda1798<=gda1798+1;	end            end
            always@(posedge clk or negedge rstn) begin	if(rstn==1'b0) begin	ribcc5<=0;	end	else begin	if(pfecd0b)	ribcc5<=ribcc5+1;	end            end
            assign mr5e62a = (gda1798 == ribcc5) ? 1'b1: 1'b0;
            always@(posedge clk or negedge rstn) begin	if(rstn==1'b0) begin	rfib<=1'b1;	end	else begin	if (((os67205)&&(!wla1295)) || mr5e62a)	rfib <= 1'b1;	else if ((ibstart&&lf94e33) || (wla1295 && !mr5e62a))	rfib <= 1'b0;	end            end  end      end      endgenerate
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module do9c345_FFTC2048 (
                clk,       
                rstn,      
                din,       
                dout       
                );
parameter fc2aae9   = 16;
input                        clk;
input                        rstn;
input  [fc2aae9-1:0]      din;
output [fc2aae9-1:0]      dout;
reg    [fc2aae9-1:0]      dout;
                              always @(posedge clk or negedge rstn) begin         if(rstn==1'b0)            dout <= 'b0;         else            dout <= din;      end
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module gdd98d_FFTC2048 (
                clk,       
                rstn,      
                ibstart,   
                dire,      
                diim,      
                ribd9a1,  
                ho5224c, 
                ph91262, 
                do89317, 
                cm498ba,     
                yk4c5d1      
                );
parameter fc2aae9   = 16;
input                        clk;
input                        rstn;
input                        ibstart;
input  [fc2aae9-1:0]      dire;
input  [fc2aae9-1:0]      diim;
output                       ribd9a1;
output                       ho5224c;
output                       ph91262;
output                       do89317;
output [fc2aae9-1:0]      cm498ba;
output [fc2aae9-1:0]      yk4c5d1;
reg                          ribd9a1;
reg                          ho5224c;
reg                          ph91262;
reg                          do89317;
reg    [fc2aae9-1:0]      cm498ba;
reg    [fc2aae9-1:0]      yk4c5d1;
                              always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ribd9a1 <= 1'b0;            ho5224c<= 1'b0;            ph91262<= 1'b0;            do89317<= 1'b0;            cm498ba <= 'b0;            yk4c5d1 <= 'b0;         end         else begin            ribd9a1 <= ibstart;            ho5224c<= ribd9a1;            ph91262<= ho5224c;            do89317<= ph91262;            cm498ba <= dire;            yk4c5d1 <= diim;         end      end
   endmodule                                                                                             
`timescale 1 ns / 100 ps
module uifa97e_FFTC2048 (
                clk,       
                rstn,      
                ibstart,   
                mode,      
                modeset,   
   
                wl80cf8      
                );
input                        clk;
input                        rstn;
input                        ibstart;
input                        mode;
input                        modeset;
output                       wl80cf8;
reg                          tu7c95b;
reg                          wl80cf8;
                           always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            tu7c95b <= 1'b0;            wl80cf8     <= 1'b0;         end         else begin            if (modeset)               tu7c95b <= mode;            if (ibstart) begin               if (modeset)                  wl80cf8 <= mode;               else                  wl80cf8 <= tu7c95b ;            end         end      end
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module ph1c7c6_FFTC2048 (
                clk,       
                rstn,      
                ibstart,   
                sfact,     
                sfactset,  
                lsbdfe5, 
                kdf8b37,
                jcc59bd,
   
                an2cdeb     
                );
parameter sfact_width   = 16;
parameter plog2_points  = 4;
parameter pdyn_points  = 0;
input                        clk;
input                        rstn;
input                        ibstart;
input  [sfact_width-1:0]     sfact;
input                        sfactset;
input  [plog2_points:0]      kdf8b37;
input                        jcc59bd;
input                        lsbdfe5;
output [sfact_width-1:0]     an2cdeb;
reg    [sfact_width-1:0]     ri9c793;
reg    [sfact_width-1:0]     ng1e4df;
reg    [sfact_width-1:0]     ls937d5;
reg    [sfact_width-1:0]     an2cdeb;
reg    [sfact_width-1:0]     fad55d0;
reg                          ho5224c;
reg                          ph91262;
wire  [plog2_points:0]	hod07d7;
reg	ri83ebb;
reg    [sfact_width-1:0]     icfaed0;
integer                      rtd7680;
genvar qvbb406;
            
                           always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ri9c793 <= {sfact_width{1'b0}};            ng1e4df  <= {sfact_width{1'b0}};         end         else begin            if (sfactset)               ri9c793 <= sfact;            if (ibstart) begin               if (sfactset)                  ng1e4df <= sfact;               else                  ng1e4df <= ri9c793 ;            end         end      end
      generate	if ((pdyn_points==1) && (plog2_points==6)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	end	else if ((pdyn_points==1) && (plog2_points==7)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	end	else if ((pdyn_points==1) && (plog2_points==8)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	end	else if ((pdyn_points==1) && (plog2_points==9)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	end	else if ((pdyn_points==1) && (plog2_points==10)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	assign hod07d7[9] = |(kdf8b37[8:0]);	end	else if ((pdyn_points==1) && (plog2_points==11)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	assign hod07d7[9] = |(kdf8b37[8:0]);	assign hod07d7[10] = |(kdf8b37[9:0]);	end	else if ((pdyn_points==1) && (plog2_points==12)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	assign hod07d7[9] = |(kdf8b37[8:0]);	assign hod07d7[10] = |(kdf8b37[9:0]);	assign hod07d7[11] = |(kdf8b37[10:0]);	end	else if ((pdyn_points==1) && (plog2_points==13)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	assign hod07d7[9] = |(kdf8b37[8:0]);	assign hod07d7[10] = |(kdf8b37[9:0]);	assign hod07d7[11] = |(kdf8b37[10:0]);	assign hod07d7[12] = |(kdf8b37[11:0]);	end	else if ((pdyn_points==1) && (plog2_points==14)) begin	assign hod07d7[2] = |(kdf8b37[1:0]);	assign hod07d7[3] = |(kdf8b37[2:0]);	assign hod07d7[4] = |(kdf8b37[3:0]);	assign hod07d7[5] = |(kdf8b37[4:0]);	assign hod07d7[6] = |(kdf8b37[5:0]);	assign hod07d7[7] = |(kdf8b37[6:0]);	assign hod07d7[8] = |(kdf8b37[7:0]);	assign hod07d7[9] = |(kdf8b37[8:0]);	assign hod07d7[10] = |(kdf8b37[9:0]);	assign hod07d7[11] = |(kdf8b37[10:0]);	assign hod07d7[12] = |(kdf8b37[11:0]);	assign hod07d7[13] = |(kdf8b37[12:0]);	end         endgenerate
      generate      begin         if (pdyn_points==1) begin
	always@(posedge clk or negedge rstn) begin	if(rstn==1'b0)	ri83ebb <= 1'b0;	else	if((ibstart)^(kdf8b37[plog2_points-1]))	ri83ebb <= ~ri83ebb;	end
                  
      always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            an2cdeb     <= {sfact_width{1'b0}};            ls937d5 <= {sfact_width{1'b0}};            icfaed0 <= {sfact_width{1'b0}};         end         else begin                                    if (ibstart)               ls937d5 <= fad55d0;                                    for (rtd7680=0;rtd7680<2;rtd7680=rtd7680+1) begin               if (kdf8b37[rtd7680]) begin                  an2cdeb[2*plog2_points-1-(2*rtd7680)]   <= fad55d0[2*plog2_points-1-(2*rtd7680)];                  an2cdeb[2*plog2_points-1-(2*rtd7680+1)] <= fad55d0[2*plog2_points-1-(2*rtd7680+1)];               end            end            for (rtd7680=2;rtd7680<plog2_points;rtd7680=rtd7680+1) begin               if (kdf8b37[rtd7680]) begin                  if ((jcc59bd&&(!hod07d7[rtd7680])) || (ri83ebb)) begin                                       an2cdeb[2*plog2_points-1-(2*rtd7680)]   <= fad55d0[2*plog2_points-1-(2*rtd7680)];
                     an2cdeb[2*plog2_points-1-(2*rtd7680+1)] <= fad55d0[2*plog2_points-1-(2*rtd7680+1)];                  end                                                                                          else begin                     an2cdeb[2*plog2_points-1-(2*rtd7680)]   <= ls937d5[2*plog2_points-1-(2*rtd7680)];                     an2cdeb[2*plog2_points-1-(2*rtd7680+1)] <= ls937d5[2*plog2_points-1-(2*rtd7680+1)];                  end               end	                                                                                                                                                   end         end      end
      always @(*) begin         if (lsbdfe5)            fad55d0 = (ng1e4df <<2);         else            fad55d0 = ng1e4df;      end
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ho5224c    <= 'b0;            ph91262    <= 'b0;         end         else begin            ho5224c    <= ibstart;            ph91262    <= ho5224c;         end      end
         end         else begin
      always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            an2cdeb     <= {sfact_width{1'b0}};            ls937d5 <= {sfact_width{1'b0}};         end         else begin            if (kdf8b37[1])               ls937d5 <= ng1e4df;            for (rtd7680=0;rtd7680<2;rtd7680=rtd7680+1) begin               if (kdf8b37[rtd7680]) begin                  an2cdeb[2*plog2_points-1-(2*rtd7680)]   <= ng1e4df[2*plog2_points-1-(2*rtd7680)];                  an2cdeb[2*plog2_points-1-(2*rtd7680+1)] <= ng1e4df[2*plog2_points-1-(2*rtd7680+1)];               end            end            for (rtd7680=2;rtd7680<plog2_points;rtd7680=rtd7680+1) begin               if (kdf8b37[rtd7680]) begin                  an2cdeb[2*plog2_points-1-(2*rtd7680)]   <= ls937d5[2*plog2_points-1-(2*rtd7680)];                  an2cdeb[2*plog2_points-1-(2*rtd7680+1)] <= ls937d5[2*plog2_points-1-(2*rtd7680+1)];               end            end         end      end
         end      end      endgenerate
   endmodule                                                                                                
`timescale 1 ns / 100 ps
module db947c_FFTC2048 (
             clk,       
             rstn,      
             ibstart,   
             points,    
             pointset,  
             kdf8b37,
             ksbc8fe,   
             mt12817,     
             lsbdfe5, 
             sw1fc5d,
             jcc59bd,
             wla1295,
             qgeff2b     
   
             );
parameter pnfft_width   = 8;
parameter plog2_points  = 4;
parameter pbfimux_level = 0;
parameter pcntmux_level = 0;
input                        clk;
input                        rstn;
input                        ibstart;
input   [pnfft_width-1:0]    points;
input                        pointset;
input   [plog2_points:0]     kdf8b37;
output  [plog2_points-1:0]   mt12817;
output                       lsbdfe5;
output  [plog2_points:0]     qgeff2b;
output  [plog2_points:0]     sw1fc5d;
output  [pnfft_width-1:0]    ksbc8fe;
output                       jcc59bd;
output                       wla1295;
reg     [pnfft_width-1:0]    ne73079;
reg     [pnfft_width-1:0]    goc1e59;
reg     [pnfft_width-1:0]    ksbc8fe;
reg     [plog2_points:0]     cm59251;
reg     [13:0]               ipc9289;
reg     [plog2_points:0]     qgeff2b;
reg     [plog2_points-1:0]   mt12817;
wire                         lsbdfe5;
wire    [pnfft_width-1:0]    ep7ac4;
wire    [pnfft_width-2:0]    xweb126;
wire    [13:0]               xw58932;
reg     [13:0]               osc4992;
reg                          ho5224c;
reg                          ph91262;
reg                          jcc59bd;
reg                          ou92227;
reg                          wla1295;
                    
                     assign sw1fc5d = osc4992;      assign xw58932  = kdf8b37;               always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ne73079 <= 'b0;            ksbc8fe     <= 'b0;            goc1e59<= 'b0;            ou92227   <= 1'b0;            wla1295  <= 1'b0;         end         else begin            ou92227     <= pointset;            if (ou92227) begin                                                                                                         goc1e59  <= ne73079;            end            if (pointset)               ne73079 <= points;            if (ibstart) begin                              if (goc1e59<6)                  ksbc8fe  <= 6;               else if (goc1e59>14)                  ksbc8fe  <= 14;               else                  ksbc8fe  <= goc1e59;            end            wla1295 <= |(ksbc8fe ^ goc1e59) ;         end      end
      assign ep7ac4 = plog2_points - ksbc8fe;      assign xweb126 = ep7ac4[pnfft_width-1:1];         generate         if (pbfimux_level==4) begin            always @(*) begin               case (xweb126)                  1: begin                     cm59251       = 4;                     osc4992[13:3] = xw58932[13:3];                     osc4992[2]    = ph91262;                     osc4992[1:0]  = xw58932[1:0];                     jcc59bd             = ph91262;                  end                  2: begin                     cm59251       = 16;                     osc4992[13:5] = xw58932[13:5];                     osc4992[4]    = ph91262;                     osc4992[3:0]  = xw58932[3:0];                     jcc59bd             = ph91262;                  end                  3: begin                     cm59251       = 64;                     osc4992[13:7] = xw58932[13:7];                     osc4992[6]    = ph91262;                     osc4992[5:0]  = xw58932[5:0];                     jcc59bd             = ph91262;                  end                  4: begin                     cm59251       = 256;                     osc4992[13:9] = xw58932[13:9];                     osc4992[8]    = ph91262;                     osc4992[7:0]  = xw58932[7:0];                     jcc59bd             = ph91262;                  end                  default: begin                     cm59251       = 0;                     osc4992[13:0] = xw58932[13:0];                     jcc59bd             = xw58932[1];                  end               endcase            end         end         if (pbfimux_level==3) begin            always @(*) begin               case (xweb126)                  1: begin                     cm59251       = 4;                     osc4992[13:3] = xw58932[13:3];                     osc4992[2]    = ph91262;                     osc4992[1:0]  = xw58932[1:0];                     jcc59bd             = ph91262;                  end                  2: begin                     cm59251       = 16;                     osc4992[13:5] = xw58932[13:5];                     osc4992[4]    = ph91262;                     osc4992[3:0]  = xw58932[3:0];                     jcc59bd             = ph91262;                  end                  3: begin                     cm59251       = 64;                     osc4992[13:7] = xw58932[13:7];                     osc4992[6]    = ph91262;                     osc4992[5:0]  = xw58932[5:0];                     jcc59bd             = ph91262;                  end                  default: begin                     cm59251       = 0;                     osc4992[13:0] = xw58932[13:0];                     jcc59bd             = xw58932[1];                  end               endcase            end         end         if (pbfimux_level==2) begin            always @(*) begin               case (xweb126)                  1: begin                     cm59251       = 4;                     osc4992[13:3] = xw58932[13:3];                     osc4992[2]    = ph91262;                     osc4992[1:0]  = xw58932[1:0];                     jcc59bd             = ph91262;                  end                  2: begin                     cm59251       = 16;                     osc4992[13:5] = xw58932[13:5];                     osc4992[4]    = ph91262;                     osc4992[3:0]  = xw58932[3:0];                     jcc59bd             = ph91262;                  end                  default: begin                     cm59251       = 0;                     osc4992[13:0] = xw58932[13:0];                     jcc59bd             = xw58932[1];                  end               endcase            end         end         if (pbfimux_level==1) begin            always @(*) begin               case (xweb126)                  1: begin                     cm59251       = 4;                     osc4992[13:3] = xw58932[13:3];                     osc4992[2]    = ph91262;                     osc4992[1:0]  = xw58932[1:0];                     jcc59bd             = ph91262;                  end                  default: begin                     cm59251       = 0;                     osc4992[13:0] = xw58932[13:0];                     jcc59bd             = xw58932[1];                  end               endcase            end         end
         if (pbfimux_level==0) begin            always @(*) begin                     cm59251       = 0;                     osc4992[13:0] = xw58932[13:0];                     jcc59bd             = xw58932[1];            end         end
      endgenerate
      
      generate         if (pcntmux_level==0) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 63;               endcase         end         if (pcntmux_level==1) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 127;               endcase         end
         if (pcntmux_level==2) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 255;               endcase         end
         if (pcntmux_level==3) begin            always @(*)               case (ksbc8fe)                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 511;               endcase         end
         if (pcntmux_level==4) begin            always @(*)               case (ksbc8fe)                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 1023;               endcase         end
         if (pcntmux_level==5) begin            always @(*)               case (ksbc8fe)                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 2047;               endcase         end
         if (pcntmux_level==6) begin            always @(*)               case (ksbc8fe)                  13:      ipc9289 = 8191;                  14:      ipc9289 = 16383;                  default: ipc9289 = 4095;               endcase         end         if (pcntmux_level==7) begin            always @(*)               case (ksbc8fe)                  14:      ipc9289 = 16383;                  default: ipc9289 = 8191;               endcase         end
         if (pcntmux_level==8) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 63;               endcase         end
         if (pcntmux_level==9) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 127;               endcase         end
         if (pcntmux_level==10) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 255;               endcase         end
         if (pcntmux_level==11) begin            always @(*)               case (ksbc8fe)                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 511;               endcase         end
         if (pcntmux_level==12) begin            always @(*)               case (ksbc8fe)                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 1023;               endcase         end
         if (pcntmux_level==13) begin            always @(*)               case (ksbc8fe)                  12:      ipc9289 = 4095;                  13:      ipc9289 = 8191;                  default: ipc9289 = 2047;               endcase         end
         if (pcntmux_level==14) begin            always @(*)               case (ksbc8fe)                  13:      ipc9289 = 8191;                  default: ipc9289 = 4095;               endcase         end
         if (pcntmux_level==15) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  default: ipc9289 = 63;               endcase         end
         if (pcntmux_level==16) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  default: ipc9289 = 127;               endcase         end
         if (pcntmux_level==17) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  default: ipc9289 = 255;               endcase         end
         if (pcntmux_level==18) begin            always @(*)               case (ksbc8fe)                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  default: ipc9289 = 511;               endcase         end
         if (pcntmux_level==19) begin            always @(*)               case (ksbc8fe)                  11:      ipc9289 = 2047;                  12:      ipc9289 = 4095;                  default: ipc9289 = 1023;               endcase         end
         if (pcntmux_level==20) begin            always @(*)               case (ksbc8fe)                  12:      ipc9289 = 4095;                  default: ipc9289 = 2047;               endcase         end
         if (pcntmux_level==21) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  default: ipc9289 = 63;               endcase         end
         if (pcntmux_level==22) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  default: ipc9289 = 127;               endcase         end         if (pcntmux_level==23) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  default: ipc9289 = 255;               endcase         end         if (pcntmux_level==24) begin            always @(*)               case (ksbc8fe)                  10:      ipc9289 = 1023;                  11:      ipc9289 = 2047;                  default: ipc9289 = 511;               endcase         end         if (pcntmux_level==25) begin            always @(*)               case (ksbc8fe)                  11:      ipc9289 = 2047;                  default: ipc9289 = 1023;               endcase         end
         if (pcntmux_level==26) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  default: ipc9289 = 63;               endcase         end
         if (pcntmux_level==27) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  default: ipc9289 = 127;               endcase         end         if (pcntmux_level==28) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  10:      ipc9289 = 1023;                  default: ipc9289 = 255;               endcase         end         if (pcntmux_level==29) begin            always @(*)               case (ksbc8fe)                  10:      ipc9289 = 1023;                  default: ipc9289 = 511;               endcase         end
         if (pcntmux_level==30) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  default: ipc9289 = 63;               endcase         end
         if (pcntmux_level==31) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  9:       ipc9289 = 511;                  default: ipc9289 = 127;               endcase         end         if (pcntmux_level==32) begin            always @(*)               case (ksbc8fe)                  9:       ipc9289 = 511;                  default: ipc9289 = 255;               endcase         end
         if (pcntmux_level==33) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  8:       ipc9289 = 255;                  default: ipc9289 = 63;               endcase         end         if (pcntmux_level==34) begin            always @(*)               case (ksbc8fe)                  8:       ipc9289 = 255;                  default: ipc9289 = 127;               endcase         end
         if (pcntmux_level==35) begin            always @(*)               case (ksbc8fe)                  7:       ipc9289 = 127;                  default: ipc9289 = 63;               endcase         end
      endgenerate
      generate         if (plog2_points%2==1)            assign lsbdfe5 = ~ksbc8fe[0];         else            assign lsbdfe5 = ksbc8fe[0];      endgenerate
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            qgeff2b    <= 'b0;            mt12817     <= 'b0;         end         else begin            qgeff2b    <= cm59251;            mt12817     <= ipc9289;         end      end
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            ho5224c    <= 'b0;            ph91262    <= 'b0;         end         else begin            ho5224c    <= ibstart;            ph91262    <= ho5224c;         end      end
   endmodule                                                                                             
`timescale 1 ns / 100 ps
module ale81d9_FFTC2048 (
            clk,       
            rstn,      
            qi5137,       
            an39028, 
            pfcdf4c, 
            os67205,  
            mt12817,     
            lsbdfe5, 
            kq4cf46,    
            kq67a31,  
            zz3d189,   
            fnc8144,      
            ip75347,       
            hd940bd,    
            ri89d08,     
            ksbc8fe,   
            except,    
            ou2b339,
            outvalid,  
            kq439ac,  
            cm599c8,  
            obstart,   
            tw35837,     
            ymac1bb  
            );
parameter pdyn_points    = 0;
parameter pnfft_width    = 8;
parameter bit_reverse    = 0;
parameter plog2_points   = 4;
parameter enc6b7b   = 16;
parameter med4d71 = "ECP";
localparam ks882e6 = 2*enc6b7b;
localparam rib864c  = (1<<plog2_points)-1;
localparam uv6579e= (1<<plog2_points)-5;
localparam kd5e7a9  = 6;
input                       clk;
input                       rstn;
input  [plog2_points:0]     qi5137;
input  [plog2_points:0]     an39028;
input  [plog2_points:0]     pfcdf4c;
input  [plog2_points+1:0]   os67205;
input  [plog2_points-1:0]   mt12817;
input                       lsbdfe5;
input                       kq4cf46;
input                       kq67a31;
input  [ks882e6-1:0]   zz3d189;
input                       fnc8144;
input                       hd940bd;
input  [ks882e6-1:0]   ri89d08;
input  [pnfft_width-1:0]    ksbc8fe;
output                      ou2b339;
output                      kq439ac;
output                      cm599c8;
output                      except;
output                      outvalid;
output                      obstart;
output                      ip75347;
output [ks882e6-1:0]   tw35837;
output   ymac1bb;
reg    [plog2_points-1:0]   hbe306d;
reg                         wl1836e;
reg                         yz7bc0;
reg    [plog2_points-1:0]   goef027;
reg                         bl6ea68;
reg                         byc09c0;
reg    [plog2_points:0]     hd2701b;
reg    [13:0]               xl380de;
reg   ymac1bb;
reg                         rv37b2;
reg                         ls1bd97;
reg                         aydecbb;
reg                         thf65d9;
reg                         zmb2ecf;
reg                         qi9767a;
reg                         irbb3d0;
reg                         uvd9e85;
reg                         rgcf42c;
reg                         qt7a163;
reg                         obstart;
reg                         outvalid;
reg                         qv2c755;
reg                         except;
reg                         yz1d56b;
reg                         ayeab5d;
reg                         bl55ae9;
reg                         riad74e;
reg                         ou2b339;
wire                        kq439ac;
wire                        cm599c8;
wire   [ks882e6-1:0]   ri89d08;
wire                        sj9f7aa;
wire                        byfbd54;
wire   [ks882e6-1:0]   tw35837;
wire                        phaa888;
wire                        qt54447;
wire                        ip75347;
wire   [plog2_points:0]     uk88f53;
wire   [plog2_points-1:0]   jp71e77;
wire   [plog2_points-1:0]   ui532b0;
wire                        fn5ff31;
wire   [ks882e6-1:0]   kq5601a;
wire                        zkc01da;
wire                        an80686;
wire   [13:0]               db3434;
integer                     rtd7680;
integer                     qvbb406;
integer                     hq869c2;
                                                      
                                 assign db3434 = goef027[plog2_points-1:0];
         generate      begin         if (pdyn_points==1) begin            assign jp71e77     = mt12817;            assign ui532b0   = mt12817 - 4;            assign fn5ff31         = lsbdfe5 ? kq67a31 :hd940bd;            assign kq5601a          = lsbdfe5 ? zz3d189  : ri89d08;            assign zkc01da = fn5ff31;            assign an80686 = qt54447;            always @(*) begin               hd2701b[plog2_points] = byc09c0;               case (ksbc8fe)                  6: begin                     xl380de[13:6] = 0;                     for(rtd7680=0;rtd7680<=5;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[5-rtd7680];                  end                  7: begin                     xl380de[13:7] = 0;                     for(rtd7680=0;rtd7680<=6;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[6-rtd7680];                  end                  8: begin                     xl380de[13:8] = 0;                     for(rtd7680=0;rtd7680<=7;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[7-rtd7680];                  end                  9: begin                     xl380de[13:9] = 0;                     for(rtd7680=0;rtd7680<=8;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[8-rtd7680];                  end                  10:begin                     xl380de[13:10] = 0;                     for(rtd7680=0;rtd7680<=9;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[9-rtd7680];                  end                  11:begin                     xl380de[13:11] = 0;                     for(rtd7680=0;rtd7680<=10;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[10-rtd7680];                  end                  12:begin                     xl380de[13:12] = 0;                     for(rtd7680=0;rtd7680<=11;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[11-rtd7680];                  end                  13:begin                     xl380de[13:13] = 0;                     for(rtd7680=0;rtd7680<=12;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[12-rtd7680];                  end                  default: begin                     for(rtd7680=0;rtd7680<=13;rtd7680=rtd7680+1)                        xl380de[rtd7680]  = db3434[13-rtd7680];                  end               endcase               hd2701b[plog2_points-1:0] = xl380de[plog2_points-1:0];            end         end         else begin            assign jp71e77     = rib864c;            assign ui532b0   = uv6579e ;            assign fn5ff31         = hd940bd ;            assign kq5601a          = ri89d08 ;            assign zkc01da = 1'b0;            assign an80686 = 1'b0;            always @(*) begin               for(rtd7680=0;rtd7680<plog2_points;rtd7680=rtd7680+1)                  hd2701b[rtd7680]=goef027[plog2_points-1-rtd7680];               hd2701b[plog2_points] = byc09c0;            end         end      end      endgenerate
         generate         if (bit_reverse==0) begin                 always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  hbe306d <= 'b0;               else if (zkc01da==1'b1)                  hbe306d <= 'b0;               else if (wl1836e==1'b1)                  hbe306d <= hbe306d+1;            end
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  wl1836e <= 1'b0;               else if (fn5ff31==1'b1)                  wl1836e <= 1'b1;               else if (phaa888==1'b1)                  wl1836e <= 1'b0;            end
               assign phaa888 = (hbe306d==jp71e77)? 1'b1 : 1'b0;
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  yz7bc0 <= 1'b0;               else if (phaa888==1'b1)                  yz7bc0 <= ~yz7bc0;            end
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  goef027 <= 'b0;               else if (an80686==1'b1)                  goef027 <= 'b0;               else if (bl6ea68==1'b1)                  goef027 <= goef027+1;            end
               assign qt54447 = (hbe306d==ui532b0)? 1'b1 : 1'b0;
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  bl6ea68 <= 1'b0;               else if (qt54447==1'b1)                  bl6ea68 <= 1'b1;               else if (ip75347==1'b1)                  bl6ea68 <= 1'b0;            end
               assign ip75347 = (goef027==jp71e77)? 1'b1 : 1'b0;
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0)                  byc09c0 <= 1'b0;               else if (qt54447==1'b1)                  byc09c0 <= yz7bc0;            end
               assign uk88f53 = {yz7bc0, hbe306d};
         
            rib7c8c_FFTC2048 #(               .ba99a50(ks882e6),               .med4d71(med4d71),               .ho69416(plog2_points+1))                    ngadc88 (                  .clk(clk),                            .rstn(rstn),                          .pfdd15f(wl1836e),                     .uk2bfe6(uk88f53),                        .neca54e(kq5601a),                      .tj9ba2b(hd2701b),                        .go7dcff(tw35837)                      );
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  rv37b2 <= 1'b0;                  ls1bd97 <= 1'b0;                  aydecbb <= 1'b0;                  thf65d9 <= 1'b0;                  zmb2ecf <= 1'b0;                  ayeab5d <= 1'b0;                  bl55ae9 <= 1'b0;                  riad74e <= 1'b0;               end               else begin                  rv37b2 <= qt54447;                  ls1bd97 <= rv37b2;                  aydecbb <= ls1bd97;                  thf65d9 <= bl6ea68;                  zmb2ecf <= thf65d9;                  ayeab5d <= ip75347;                  bl55ae9 <= ayeab5d;                  riad74e <= bl55ae9;               end            end
               assign kq439ac  = ls1bd97;            assign sj9f7aa = zmb2ecf;            assign byfbd54= thf65d9;            assign cm599c8 = aydecbb;
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  yz1d56b   <= 1'b0;               end               else begin                  if (aydecbb)                     yz1d56b   <= 1'b0 ;                  for(hq869c2=1;hq869c2<plog2_points;hq869c2=hq869c2+1) begin                     if (os67205[hq869c2])                        yz1d56b   <= yz1d56b | pfcdf4c[hq869c2];                     if (ls1bd97)                        yz1d56b   <= yz1d56b | pfcdf4c[plog2_points];                  end               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  except   <= 1'b0;               end               else begin                  if ((yz1d56b)&&(cm599c8))                     except   <= 1'b1;                  else if (riad74e)                     except   <= 1'b0;               end            end
         end         else begin               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  uvd9e85     <= 1'b0;                  rgcf42c   <= 1'b0;                  qt7a163     <= 1'b0;                  qi9767a   <= 1'b0;                  irbb3d0 <= 1'b0;                  qv2c755  <= 1'b0;               end               else begin                  uvd9e85     <= fnc8144;                  rgcf42c   <= kq4cf46;                  qt7a163     <= uvd9e85;                  qi9767a   <= hd940bd;                  irbb3d0 <= kq67a31;                  qv2c755  <= fn5ff31;               end            end            assign kq439ac  = fn5ff31;            assign sj9f7aa = lsbdfe5 ? rgcf42c     : uvd9e85;            assign byfbd54= lsbdfe5 ? kq4cf46        : fnc8144;            assign cm599c8  = qv2c755;            assign tw35837    = kq5601a;
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                                    ou2b339   <= 1'b0;               end               else begin                  if (cm599c8)                     ou2b339   <= ~ou2b339;               end            end
               always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  yz1d56b   <= 1'b0;               end               else begin                                                                                                                                                                  yz1d56b   <= |pfcdf4c[plog2_points:1];               end            end
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  except   <= 1'b0;               end               else begin                  if (cm599c8)                     except   <= yz1d56b;                  else if (sj9f7aa) begin                     if ((yz1d56b)||(except))                     except   <= 1'b1;                  end                  else                     except   <= 1'b0;               end            end
         end      endgenerate
         always @(posedge clk or negedge rstn) begin         if(rstn==1'b0) begin            outvalid   <= 1'b0;            obstart    <= 1'b0;         end         else begin            outvalid   <= sj9f7aa;            ymac1bb <= byfbd54;            obstart    <= cm599c8;         end      end
   endmodule                                                                                    
`timescale 1 ns / 100 ps
module yzb4add_FFTC2048 (
            clk,                  
            rstn,                 
            din,                  
            cz709f8,                
            qgeff2b,               
            except,               
            dout                  
          ) ;
parameter pdyn_points    = 0;
parameter twb8d6f    = 0;
parameter fc2aae9     = 16;
parameter epaba5f    = 16;
parameter fixed_scaling  = 1;
parameter rounding_method= 1;
parameter pscale_reg     = 0;
parameter plog2_points   = 4;
parameter ptrunc_laststgs= 0;
input                      clk;
input                      rstn;
input [fc2aae9-1:0]     din;
input [1:0]                cz709f8;
input                      qgeff2b;
output                     except;
output [epaba5f-1:0]   dout;
reg  [epaba5f-1:0]     yz9a957;
wire [epaba5f-1:0]     dout;
wire                       except;
wire                       ne57a3b;
reg  [fc2aae9-1:0]      ene8eda;
reg                        by476d4;
reg                        mg3b6a3;
wire                       ykdb519;
                                                
   
                           assign ne57a3b = din[fc2aae9-1] ;      assign except = 1'b0;
                     generate         if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-1:1];         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-1:1];                  end                  2'b10 : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-1:2]};                  end                  default : begin                     yz9a957 = din[fc2aae9-2:0];                  end               endcase            end            assign dout = yz9a957;         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-1:1];         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-1:1];                  end                  2'b10 : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-1:2]};                  end                  default : begin                     yz9a957 = din[fc2aae9-2:0];                  end               endcase            end            assign dout = yz9a957;         end         else if ((fixed_scaling==3) && (rounding_method==1)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = ene8eda[fc2aae9-1:1];                  end                  2'b10 : begin                     yz9a957 = {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]};                  end                  default : begin                     yz9a957 = ene8eda[fc2aae9-2:0];                  end               endcase            end            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;               end               else begin                  ene8eda  <= din;               end            end            assign dout = yz9a957;         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-1:1];         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]);                  end                  2'b10 : begin                     yz9a957 = ne57a3b ? ({din[fc2aae9-1],din[fc2aae9-1:2]}+(din[1]&din[0]))                                 : {din[fc2aae9-1],din[fc2aae9-1:2]}+din[1];                  end                  default : begin                     yz9a957 = din[fc2aae9-1:0];                  end               endcase            end            assign dout = yz9a957;         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-1:1];         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]);                  end                  2'b10 : begin                     yz9a957 = ne57a3b ? ({din[fc2aae9-1],din[fc2aae9-1:2]}+(din[1]&din[0]))                                 : {din[fc2aae9-1],din[fc2aae9-1:2]}+din[1];                  end                  default : begin                     yz9a957 = din[fc2aae9-1:0];                  end               endcase            end            assign dout = yz9a957;         end         else if ((fixed_scaling==3) && (rounding_method==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0]);                  end                  2'b10 : begin                     yz9a957 = by476d4 ? ({ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+(ene8eda[1]&ene8eda[0]))                                 : {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+ene8eda[1];                  end                  default : begin                     yz9a957 = ene8eda[fc2aae9-1:0];                  end               endcase            end            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout = yz9a957;         end                  else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==1)&&(pdyn_points==0)) begin            assign dout[epaba5f-1:0] = {din[fc2aae9-1],din[fc2aae9-1:2]};         end         else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==1)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;               end               else begin                  ene8eda  <= din;               end            end            assign dout[epaba5f-1:0] = {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}  ;         end         else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = by476d4 ? ({ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+(ene8eda[1]&ene8eda[0]))                                              : {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+ene8eda[1]  ;         end         else if  ((fixed_scaling==2) && (rounding_method==1)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1];         end         else if  ((fixed_scaling==2) && (rounding_method==1)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  mg3b6a3   <= 1'b0;               end               else begin                  ene8eda  <= din;                  mg3b6a3   <= qgeff2b;               end            end            assign dout[epaba5f-1:0] = mg3b6a3 ? {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]} : ene8eda[fc2aae9-1:1]  ;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = qgeff2b ? (ne57a3b ? ({din[fc2aae9-1],din[fc2aae9-1:2]}+(din[1]&din[0])) : {din[fc2aae9-1],din[fc2aae9-1:2]}+din[1] ) : (ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ) ;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;                  mg3b6a3   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= 
ne57a3b;                  mg3b6a3   <= qgeff2b;               end            end            assign dout[epaba5f-1:0] = mg3b6a3 ? (by476d4 ? ({ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+(ene8eda[1]&ene8eda[0])) : {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+ene8eda[1] ) : (by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0]) )  ;         end
         else if  ((fixed_scaling==2) && (rounding_method==1)&&(pdyn_points==0)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1];         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(pdyn_points==0)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(pdyn_points==0)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(pdyn_points==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0])  ;         end
                  else if  ((fixed_scaling==1) && (rounding_method==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ;         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ;         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f!=(plog2_points-1))) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0])  ;         end
      endgenerate
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module pua7955_FFTC2048 (
            clk,                  
            rstn,                 
            din,                  
            cz709f8,                
            qgeff2b,               
            except,               
            dout                  
          ) ;
parameter pdyn_points    = 0;
parameter twb8d6f    = 0;
parameter fc2aae9     = 16;
parameter epaba5f    = 16;
parameter fixed_scaling  = 1;
parameter rounding_method= 1;
parameter pscale_reg     = 0;
parameter plog2_points   = 4;
parameter ptrunc_laststgs= 0;
input                      clk;
input                      rstn;
input [fc2aae9-1:0]     din;
input [1:0]                cz709f8;
input                      qgeff2b;
output                     except;
output [epaba5f-1:0]   dout;
reg  [epaba5f-1:0]     yz9a957;
wire [epaba5f-1:0]     dout;
wire                       except;
wire                       ne57a3b;
reg  [fc2aae9-1:0]      ene8eda;
reg                        by476d4;
reg                        mg3b6a3;
reg                        ykdb519;
reg [fc2aae9-1:0]    aa3eb56;
reg [fc2aae9-1:0]    twad581;
                                                
   
                     always @(posedge clk or negedge rstn) begin            if(!rstn) begin               aa3eb56   <= 0;               twad581 <= 0;            end            else begin               aa3eb56   <= din;               twad581 <= ene8eda;            end         end
         assign ne57a3b = din[fc2aae9-1] ;
                     generate         if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-2:0];            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-2:0];                     ykdb519 = ^aa3eb56[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = din[fc2aae9-1:1];                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-3:0],1'b0};                     ykdb519 = (|aa3eb56[fc2aae9-1:fc2aae9-3])&(!(&aa3eb56[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            assign dout = yz9a957;            assign except = ykdb519;         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-2:0];            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if ((fixed_scaling==3) && (rounding_method==1)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-2:0];                     ykdb519 = ^aa3eb56[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = din[fc2aae9-1:1];                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-3:0],1'b0};                     ykdb519 = (|aa3eb56[fc2aae9-1:fc2aae9-3])&(!(&aa3eb56[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            assign dout = yz9a957;            assign except = ykdb519;         end         else if ((fixed_scaling==3) && (rounding_method==1)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = ene8eda[fc2aae9-2:0];                     ykdb519 = ^twad581[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = ene8eda[fc2aae9-1:1];                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {ene8eda[fc2aae9-1],ene8eda[fc2aae9-3:0],1'b0};                     ykdb519 = (|twad581[fc2aae9-1:fc2aae9-3])&(!(&twad581[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;               end               else begin                  ene8eda  <= din;               end            end            assign dout = yz9a957;            assign except = ykdb519;         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-2:0];            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-2:0] ;                     ykdb519 = ^aa3eb56[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]);                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-3:0],1'b0};                     ykdb519 = (|aa3eb56[fc2aae9-1:fc2aae9-3])&(!(&aa3eb56[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            assign dout = yz9a957;            assign except = ykdb519;         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout = din[fc2aae9-2:0];            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if ((fixed_scaling==3) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = din[fc2aae9-2:0] ;                     ykdb519 = ^aa3eb56[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]);                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {din[fc2aae9-1],din[fc2aae9-3:0],1'b0};                     ykdb519 = (|aa3eb56[fc2aae9-1:fc2aae9-3])&(!(&aa3eb56[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            assign dout = yz9a957;            assign except = ykdb519;         end         else if ((fixed_scaling==3) && (rounding_method==0)) begin            always @(*) begin               case (cz709f8)                  2'b01 : begin                     yz9a957 = ene8eda[fc2aae9-2:0] ;                     ykdb519 = ^twad581[fc2aae9-1:fc2aae9-2];                  end                  2'b10 : begin                     yz9a957 = by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0]);                     ykdb519 = 1'b0;                  end                  default : begin                     yz9a957 = {ene8eda[fc2aae9-1],ene8eda[fc2aae9-3:0],1'b0};                     ykdb519 = (|twad581[fc2aae9-1:fc2aae9-3])&(!(&twad581[fc2aae9-1:fc2aae9-3]));                  end               endcase            end            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout = yz9a957;            assign except = ykdb519;         end                  else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==1)&&(pdyn_points==0)) begin            assign dout[epaba5f-1:0] = {din[fc2aae9-1],din[fc2aae9-1:2]};            assign except = 1'b0;         end         else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==1)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;               end               else begin                  ene8eda  <= din;               end            end            assign dout[epaba5f-1:0] = {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}  ;            assign except = 1'b0;         end         else if ((fixed_scaling==2) && (twb8d6f==0) && (rounding_method==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = by476d4 ? ({ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+(ene8eda[1]&ene8eda[0]))                                              : {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+ene8eda[1]  ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==1)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1];            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==1)&&(pdyn_points==1)) begin
            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  mg3b6a3   <= 1'b0;               end               else begin                  ene8eda  <= din;                  mg3b6a3   <= qgeff2b;               end            end            assign dout[epaba5f-1:0] = mg3b6a3 ? {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]} : ene8eda[fc2aae9-1:1]  ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&((twb8d6f==(plog2_points-1))||(twb8d6f==(plog2_points-2)))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = qgeff2b ? (ne57a3b ? ({din[fc2aae9-1],din[fc2aae9-1:2]}+(din[1]&din[0])) : {din[fc2aae9-1],din[fc2aae9-1:2]}+din[1] ) : (ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ) ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(pdyn_points==1)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;                  mg3b6a3   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;                  mg3b6a3   <= qgeff2b;               end            end            assign dout[epaba5f-1:0] = mg3b6a3 ? (by476d4 ? ({ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+(ene8eda[1]&ene8eda[0])) : {ene8eda[fc2aae9-1],ene8eda[fc2aae9-1:2]}+ene8eda[1] ) : (by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0]) )  ;            assign except = 1'b0;         end
         else if  ((fixed_scaling==2) && (rounding_method==1)&&(pdyn_points==0)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1];            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(pdyn_points==0)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-1:1] ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(pdyn_points==0)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = ne57a3b ? din[fc2aae9-1:1] : (din[fc2aae9-1:1]+din[0]) ;            assign except = 1'b0;         end         else if  ((fixed_scaling==2) && (rounding_method==0)&&(pdyn_points==0)) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = by476d4 ? ene8eda[fc2aae9-1:1] : (ene8eda[fc2aae9-1:1]+ene8eda[0])  ;            assign except = 1'b0;         end
                  else if  ((fixed_scaling==1) && (rounding_method==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-2:0];            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-2:0] ;            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-1))&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-2:0] ;            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==1)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-2:0] ;            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f==(plog2_points-2))&&(pdyn_points==1)&&(ptrunc_laststgs==0)) begin            assign dout[epaba5f-1:0] = din[fc2aae9-2:0] ;            assign except = ^aa3eb56[fc2aae9-1:fc2aae9-2];         end         else if  ((fixed_scaling==1) && (rounding_method==0)&&(twb8d6f!=(plog2_points-1))) begin            always @(posedge clk or negedge rstn) begin               if(rstn==1'b0) begin                  ene8eda  <= 'b0;                  by476d4   <= 1'b0;               end               else begin                  ene8eda  <= din;                  by476d4   <= ne57a3b;               end            end            assign dout[epaba5f-1:0] = ene8eda[fc2aae9-2:0] ;            assign except = ^twad581[fc2aae9-1:fc2aae9-2];         end
      endgenerate
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module ofdc411_FFTC2048 (
            clk,      
            rstn,     
            ks82361,    
            hq11b09,    
            mg8d84a      
            );
parameter by6c251 = 16;
parameter jp6128b = 16;
parameter rv945f=0;
parameter device_family = "ECP2";
localparam kd517f7=by6c251+jp6128b;
input                       clk;
input                       rstn;
input  [by6c251-1:0]    ks82361;
input  [jp6128b-1:0]    hq11b09;
output [kd517f7-1:0]     mg8d84a;
wire   [by6c251-1:0]    ks82361;
wire   [jp6128b-1:0]    hq11b09;
wire   [kd517f7-1:0]     mg8d84a;
                                                                                             pmi_mult #( .pmi_dataa_width           (by6c251   ),                         .pmi_datab_width           (jp6128b   ),                         .module_type               ("pmi_mult"    ),                         .pmi_sign                  ("on"          ),                         .pmi_additional_pipeline   (rv945f),                         .pmi_input_reg             ("off"          ),                         .pmi_output_reg            ("off"          ),                         .pmi_family                (device_family ),                         .pmi_implementation        ("LUT"         ))         ie8271c (                     .DataA                     (ks82361         ),                     .DataB                     (hq11b09         ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (mg8d84a          )                  );
   endmodule                                                                                             
`timescale 1 ns / 100 ps
module tue1eff_FFTC2048 (
               clk,              
               rstn,             
               bydfe8e,
               dout              
               );
parameter qgfa399    = 10;
parameter ead1cc9    = 16;
parameter rv8e648    = "reg";
parameter ps73247  = "twidFFTC2048.mem";
parameter tw9923b     = "ECP2";
parameter ofc91db    = 1;
parameter ne48edc     = 1024;
parameter jc476e3 = qgfa399-2;
parameter qgdb8d9     = 1<<qgfa399;
parameter rte364d    = qgdb8d9/4;
parameter qtd9372    = qgdb8d9/2;
parameter ho4dcad = 1<<jc476e3;
parameter kq72b5e    = ho4dcad * ead1cc9;
input                      clk;
input                      rstn;
input [qgfa399-1:0] bydfe8e;
output[ead1cc9*2-1:0] dout;
reg [ead1cc9-1:0]   dme1d4e ;
reg [ead1cc9-1:0]   wj75392 ;
reg [qgfa399-3:0]   kd4e4a0;
reg [qgfa399-3:0]   ec92829;
reg [1:0]               vx94149;
reg [1:0]               bna0a4f;
wire[ead1cc9-1:0]   mt293f0;
wire[ead1cc9-1:0]   jp4fc29;
wire[1:0]                  bl7e14e;
wire[1:0]                  osf0a77;
reg [1:0]   mt853b9;
reg [1:0]   ux29dcc;
wire[ead1cc9-1:0]   ea77324;
wire[ead1cc9-1:0]   uvcc909;
reg [ead1cc9-1:0]   gq2426e;
reg [ead1cc9-1:0]   vx9b89;
reg [1:0]   vi4dc4f;
reg [1:0]   xj6e27b;
wire[ead1cc9-1:0]   ri89ef6 = {1'b0,{(ead1cc9-1){1'b1}}};
wire[ead1cc9-1:0]   icdecfe = {1'b1,{(ead1cc9-2){1'b0}},1'b1};
assign dout = {dme1d4e,wj75392};
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            kd4e4a0 <= 0;         else if(bydfe8e[qgfa399-2])            kd4e4a0 <= -{1'b0, bydfe8e[qgfa399-3:0]};         else            kd4e4a0 <= bydfe8e[qgfa399-3:0];      end      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ec92829 <= 0;         else if(bydfe8e[qgfa399-2])            ec92829 <= bydfe8e[qgfa399-3:0];         else            ec92829 <= -{1'b0, bydfe8e[qgfa399-3:0]};      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            vx94149 <= 2'b00;         else if(bydfe8e==rte364d)            vx94149 <= 2'b01;         else if(bydfe8e>qtd9372)            vx94149 <= 2'b10;         else            vx94149 <= 2'b11;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            bna0a4f <= 2'b00;         else if(bydfe8e==0)            bna0a4f <= 2'b01;         else if(bydfe8e==qtd9372)            bna0a4f <= 2'b10;         else if(bydfe8e<=rte364d)            bna0a4f <= 2'b11;         else            bna0a4f <= 2'b00;      end
      generate      begin         if((ofc91db==0)||((ofc91db==2)&&(kq72b5e>ne48edc))) begin              pmi_ram_dp_true #(.pmi_addr_depth_a (ho4dcad   ),                              .pmi_addr_width_a (jc476e3   ),                              .pmi_data_width_a (ead1cc9   ),                              .pmi_addr_depth_b (ho4dcad   ),                              .pmi_addr_width_b (jc476e3   ),                              .pmi_data_width_b (ead1cc9   ),                              .pmi_regmode_a    (rv8e648      ),                              .pmi_regmode_b    (rv8e648      ),                              .pmi_init_file    (ps73247    ),                              .pmi_init_file_format ("binary"      ),                              .pmi_gsr          ("disable"          ),                              .pmi_resetmode    ("sync"            ),                              .pmi_write_mode_a ("normal"          ),                              .pmi_write_mode_b ("normal"          ),                              .pmi_family       (tw9923b       ),                              .module_type      ("pmi_ram_dp_true"))            dm47c23 (                              .DataInA    (           ),                              .DataInB    (           ),                              .AddressA   (ec92829    ),                              .AddressB   (kd4e4a0    ),                              .ClockA     (clk        ),                              .ClockB     (clk        ),                              .ClockEnA   (1'b1       ),                              .ClockEnB   (1'b1       ),                              .WrA        (1'b0       ),                              .WrB        (1'b0       ),                              .ResetA     (1'b0       ),                              .ResetB     (1'b0       ),                              .QA         (mt293f0  ),                              .QB         (jp4fc29  )                           );
         end else begin                pmi_distributed_rom   #(.pmi_addr_depth   (ho4dcad       ),                                    .pmi_addr_width   (jc476e3       ),                                    .pmi_data_width   (ead1cc9       ),                                    .pmi_regmode      (rv8e648          ),                                    .pmi_init_file    (ps73247        ),                                    .pmi_init_file_format ("binary"          ),                                    .pmi_family       (tw9923b           ),                                    .module_type      ("pmi_distributed_rom"))            qg5cdd2 (                                    .Address          (ec92829    ),                                    .OutClock         (clk        ),                                    .OutClockEn       (1'b1       ),                                    .Reset            (1'b0       ),                                    .Q                (ea77324  )                                    );            pmi_distributed_rom   #(.pmi_addr_depth   (ho4dcad       ),                                    .pmi_addr_width   (jc476e3       ),                                    .pmi_data_width   (ead1cc9       ),                                    .pmi_regmode      (rv8e648          ),                                    .pmi_init_file    (ps73247        ),                                    .pmi_init_file_format ("binary"          ),                                    .pmi_family       (tw9923b           ),                                    .module_type      ("pmi_distributed_rom"))            byf4082 (                                    .Address          (kd4e4a0    ),                                    .OutClock         (clk        ),                                    .OutClockEn       (1'b1       ),                                    .Reset            (1'b0       ),                                    .Q                (uvcc909  )                                    );
            always @(posedge clk or negedge rstn)            begin               if(!rstn) begin                  gq2426e <= 0;                  vx9b89 <= 0;               end else begin                  gq2426e <= ea77324;                  vx9b89 <= uvcc909;               end            end            assign mt293f0 = gq2426e;            assign jp4fc29 = vx9b89;         end         if(rv8e648=="reg") begin            always @(posedge clk or negedge rstn)            begin               if(!rstn) begin                  vi4dc4f <= 2'b00;                  xj6e27b <= 2'b00;                  mt853b9  <= 2'b00;                  ux29dcc  <= 2'b00;               end else begin                  vi4dc4f <= vx94149;                  xj6e27b <= bna0a4f;                  mt853b9  <= vi4dc4f;                  ux29dcc  <= xj6e27b;               end            end         end else begin            always @(posedge clk or negedge rstn)            begin               if(!rstn) begin                  mt853b9  <= 2'b00;                  ux29dcc  <= 2'b00;               end else begin                  mt853b9  <= vx94149;                  ux29dcc  <= bna0a4f;               end            end         end         assign bl7e14e = mt853b9;         assign osf0a77 = ux29dcc;      end      endgenerate
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            dme1d4e <= 0;         else case(osf0a77)            2'b00 : dme1d4e <= 0 - mt293f0;            2'b01 : dme1d4e <= ri89ef6;            2'b10 : dme1d4e <= icdecfe;            2'b11 : dme1d4e <= mt293f0;         endcase      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            wj75392 <= 0;         else case(bl7e14e)            2'b00 : wj75392 <= 0;            2'b01 : wj75392 <= icdecfe;            2'b10 : wj75392 <= jp4fc29;            2'b11 : wj75392 <= 0 - jp4fc29;         endcase      end
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module osf5e4e_FFTC2048 (
            clk,       
            rstn,      
            ph38443,    
            ri110f7,    
            wlbe0cb,    
            zm832e8,    
            hbd80ed,   
            ph3b7a    
            );
parameter pdin_widthr     = 16;
parameter xj71cad     = 16;
parameter phard_mac       = 1;
parameter sw31626      = 0;
parameter ph8b130= 1;
parameter zk58987  = 0;
parameter plog2_points    = 10;
parameter hqadee3      = 1;
parameter xyadfc4   = 16;
parameter device_family   = "ECP2";
input                       clk;
input                       rstn;
input  [pdin_widthr-1:0]    ph38443;
input  [pdin_widthr-1:0]    ri110f7;
input  [xj71cad-1:0]    wlbe0cb;
input  [xj71cad-1:0]    zm832e8;
output [pdin_widthr-1:0]    hbd80ed;
output [pdin_widthr-1:0]    ph3b7a;
wire                        clk;
wire                        rstn;
wire   [pdin_widthr-1:0]    ph38443;
wire   [pdin_widthr-1:0]    ri110f7;
wire   [xj71cad-1:0]    wlbe0cb;
wire   [xj71cad-1:0]    zm832e8;
wire   [pdin_widthr-1:0]    hbd80ed;
wire   [pdin_widthr-1:0]    ph3b7a;
                                                            
                           generate         if(phard_mac==1)            uieff46_FFTC2048 # (               .hqadee3(hqadee3),               .pdin_widthr(pdin_widthr),               .xj71cad(xj71cad),               .plog2_points (plog2_points),               .xyadfc4(xyadfc4),               .device_family(device_family)               )            zkf13a4 (               .clk(clk),                         .rstn(rstn),                       .ph38443(ph38443),                   .ri110f7(ri110f7),                   .wlbe0cb(wlbe0cb),                   .zm832e8(zm832e8),                   .hbd80ed(hbd80ed),                 .ph3b7a(ph3b7a)                  );
         else            ayce5bc_FFTC2048 # (               .hqadee3(hqadee3),               .pdin_widthr(pdin_widthr),               .xj71cad(xj71cad),               .device_family(device_family)               )            lqd0708 (               .clk(clk),                         .rstn(rstn),                       .ph38443(ph38443),                   .ri110f7(ri110f7),                   .wlbe0cb(wlbe0cb),                   .zm832e8(zm832e8),                   .hbd80ed(hbd80ed),                 .ph3b7a(ph3b7a)                  );
      endgenerate
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module rib7c8c_FFTC2048 (
            clk,       
            rstn,      
            pfdd15f,     
            uk2bfe6,     
            neca54e,    
            tj9ba2b,     
            go7dcff    
            );
parameter ba99a50      = 16;
parameter ho69416      = 16;
parameter gq1a9ae     = 1;
parameter med4d71 = "ECP";
localparam kqde610   = 1<<ho69416;
input                      clk;
input                      rstn;
input                      pfdd15f;
input  [ho69416-1:0]     uk2bfe6;
input  [ba99a50-1:0]     neca54e;
input  [ho69416-1:0]     tj9ba2b;
output [ba99a50-1:0]     go7dcff;
reg    [ba99a50-1:0]     uv5be0e;
wire   [ba99a50-1:0]     alf83aa;
wire                       cmc1d54;
wire                       vkeaa1;
reg    [ba99a50-1:0]     phaa854;
                                          assign cmc1d54 = 1'b1;      assign vkeaa1 = 1'b1;
      generate
      if (gq1a9ae==0) begin         pmi_distributed_dpram  #(            .pmi_addr_depth (kqde610),            .pmi_addr_width (ho69416),            .pmi_data_width (ba99a50),            .pmi_regmode    ("reg"),            .pmi_init_file  ("none"),            .pmi_init_file_format ("binary"),            .module_type    ("pmi_distributed_dpram"),            .pmi_family     (med4d71)            )            ea688fd (               .WrAddress   (uk2bfe6),               .Data        (neca54e),               .WrClock     (clk),               .WE          (pfdd15f),               .WrClockEn   (vkeaa1),               .RdAddress   (tj9ba2b),               .RdClock     (clk),               .RdClockEn   (cmc1d54),               .Reset       (~rstn),               .Q           (alf83aa)               );
         assign go7dcff = alf83aa;
      end      else         pmi_ram_dp #(            .pmi_wr_addr_depth (kqde610),            .pmi_wr_addr_width (ho69416),            .pmi_wr_data_width (ba99a50),            .pmi_rd_addr_depth (kqde610),            .pmi_rd_addr_width (ho69416),            .pmi_rd_data_width (ba99a50),            .pmi_regmode       ("reg"),            .pmi_gsr           ("disable"),            .pmi_init_file     ("none"),            .pmi_init_file_format ("binary"),            .pmi_resetmode     ("sync"),            .module_type       ("pmi_ram_dp"),            .pmi_family        (med4d71)            )         ui536e7 (               .WrAddress   (uk2bfe6),               .RdAddress   (tj9ba2b),               .Data        (neca54e),               .RdClock     (clk),               .WrClock     (clk),               .RdClockEn   (cmc1d54),               .WrClockEn   (vkeaa1),               .WE          (pfdd15f),               .Reset       (1'b0),               .Q           (go7dcff)               );
      endgenerate
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module uieff46_FFTC2048 (
            clk,       
            rstn,      
            ph38443,    
            ri110f7,    
            wlbe0cb,    
            zm832e8,    
            hbd80ed,   
            ph3b7a    
            );
parameter pdin_widthr     = 16;
parameter xj71cad     = 16;
parameter sw31626      = 0;
parameter ph8b130= 1;
parameter zk58987  = 0;
parameter plog2_points    = 10;
parameter hqadee3      = 1;
parameter xyadfc4   = 16;
parameter device_family   = "ECP2";
localparam blc24ca = pdin_widthr+xj71cad;
localparam pu995e2 = pdin_widthr+xj71cad+1;
localparam gqbc4d3 = (hqadee3==2)? (blc24ca-2) : (blc24ca-1);
localparam kdd3134   = (hqadee3==2)? (xj71cad-1): xj71cad;
localparam pf611f7 = xyadfc4+plog2_points;
localparam ie3efea = (xyadfc4==pdin_widthr)?pdin_widthr:pf611f7;
localparam kd5b896 = ie3efea + xj71cad +1;
localparam mt12d6c = ie3efea-pdin_widthr;
localparam baad95f = device_family=="ECP3" ? "on" : "off";
input                       clk;
input                       rstn;
input  [pdin_widthr-1:0]    ph38443;
input  [pdin_widthr-1:0]    ri110f7;
input  [xj71cad-1:0]    wlbe0cb;
input  [xj71cad-1:0]    zm832e8;
output [pdin_widthr-1:0]    hbd80ed;
output [pdin_widthr-1:0]    ph3b7a;
wire   [pdin_widthr-1:0]    ph38443;
wire   [pdin_widthr-1:0]    ri110f7;
wire   [xj71cad-1:0]    wlbe0cb;
wire   [xj71cad-1:0]    zm832e8;
wire   [pdin_widthr-1:0]    hbd80ed;
wire   [pdin_widthr-1:0]    ph3b7a;
reg    [ie3efea-1:0]     hbd2544;
reg    [ie3efea-1:0]     gd95131;
wire   [kd5b896-1:0]     qt44c6a;
wire   [kd5b896-1:0]     wy31aac;
integer                     rtd7680,qvbb406;
                                                                              
      
            
      
                                          always @(ph38443) begin         for(rtd7680=0;rtd7680<mt12d6c;rtd7680=rtd7680+1)            hbd2544[ie3efea-1-rtd7680]=ph38443[pdin_widthr-1];         hbd2544[pdin_widthr-1:0]=ph38443;      end
      always @(ri110f7) begin         for(qvbb406=0;qvbb406<mt12d6c;qvbb406=qvbb406+1)            gd95131[ie3efea-1-qvbb406]=ri110f7[pdin_widthr-1];         gd95131[pdin_widthr-1:0]=ri110f7;      end
                  pmi_dsp_multaddsub #( .pmi_dataa_width        (ie3efea       ),                               .pmi_datab_width        (xj71cad      ),                               .module_type            ("pmi_dsp_multaddsub" ),                               .pmi_additional_pipeline(1                ),                               .pmi_input_reg          ("on"             ),                               .pmi_output_reg         ("on"             ),                               .pmi_family             (device_family    ),                               .pmi_pipelined_mode     (baad95f    ))         bnba6f5 (.A0           (hbd2544         ),                     .A1           (gd95131         ),                     .B0           (wlbe0cb         ),                     .B1           (zm832e8         ),                     .SRIA         (               ),                     .SRIB         (               ),                     .CLK0         (clk            ),                     .CLK1         (clk            ),                     .CLK2         (clk            ),                     .CLK3         (clk            ),                     .CE0          (1'b1           ),                     .CE1          (1'b1           ),                     .CE2          (1'b1           ),                     .CE3          (1'b1           ),                     .RST0         (1'b0           ),                     .RST1         (1'b0           ),                     .RST2         (1'b0           ),                     .RST3         (1'b0           ),                     .SignA        (1'b1           ),                     .SignB        (1'b1           ),                     .ShiftA0      (1'b0           ),                     .ShiftA1      (1'b0           ),                     .ShiftB0      (1'b0           ),                     .ShiftB1      (1'b0           ),                     .ADDNSUB      (1'b0           ),                     .SUM          (qt44c6a         ),                     .SROA         (               ),                     .SROB         (               ));                  pmi_dsp_multaddsub #( .pmi_dataa_width        (ie3efea       ),                               .pmi_datab_width        (xj71cad      ),                               .module_type            ("pmi_dsp_multaddsub" ),                               .pmi_additional_pipeline(1                ),                               .pmi_input_reg          ("on"             ),                               .pmi_output_reg         ("on"             ),                               .pmi_family             (device_family    ),                               .pmi_pipelined_mode     (baad95f    ))         ls25fa2 (.A0           (hbd2544         ),                     .A1           (gd95131         ),                     .B0           (zm832e8         ),                     .B1           (wlbe0cb         ),                     .SRIA         (               ),                     .SRIB         (               ),                     .CLK0         (clk            ),                     .CLK1         (clk            ),                     .CLK2         (clk            ),                     .CLK3         (clk            ),                     .CE0          (1'b1           ),                     .CE1          (1'b1           ),                     .CE2          (1'b1           ),                     .CE3          (1'b1           ),                     .RST0         (1'b0           ),                     .RST1         (1'b0           ),                     .RST2         (1'b0           ),                     .RST3         (1'b0           ),                     .SignA        (1'b1           ),                     .SignB        (1'b1           ),                     .ShiftA0      (1'b0           ),                     .ShiftA1      (1'b0           ),                     .ShiftB0      (1'b0           ),                     .ShiftB1      (1'b0           ),                     .ADDNSUB      (1'b1           ),                     .SUM          (wy31aac         ),                     .SROA         (               ),                     .SROB         (               ));                                                                                                                                                                                             
         assign hbd80ed = qt44c6a[gqbc4d3:kdd3134];      assign ph3b7a = wy31aac[gqbc4d3:kdd3134];
   endmodule                                                                                                         
`timescale 1 ns / 100 ps
module ayce5bc_FFTC2048 (
            clk,       
            rstn,      
            ph38443,    
            ri110f7,    
            wlbe0cb,    
            zm832e8,    
            hbd80ed,   
            ph3b7a    
            );
parameter pdin_widthr   = 16;
parameter xj71cad   = 16;
parameter ui7de82 = 1;
parameter kqef411 = 1;
parameter yx7a088   = 1;
parameter hqadee3      = 1;
parameter device_family   = "ECP2";
localparam blc24ca = pdin_widthr+xj71cad;
localparam co2b2ce = pdin_widthr*2;
localparam gqbc4d3 = (hqadee3==2)? (blc24ca-2) : (blc24ca-1);
localparam kdd3134   = (hqadee3==2)? (xj71cad-1): xj71cad;
input                                       clk;
input                                       rstn;
input  [pdin_widthr-1:0]    ph38443;
input  [pdin_widthr-1:0]    ri110f7;
input  [xj71cad-1:0]    wlbe0cb;
input  [xj71cad-1:0]    zm832e8;
output [pdin_widthr-1:0]    hbd80ed;
output [pdin_widthr-1:0]    ph3b7a;
reg    [co2b2ce-1:0]   en44dc6;
wire   [blc24ca-1:0]     xw63336;
wire   [blc24ca-1:0]     alccd96;
wire   [blc24ca-1:0]     qv365ab;
wire   [blc24ca-1:0]     hq96aea;
wire   [blc24ca-1:0]     wlaba9e;
wire   [blc24ca-1:0]     meea7ab;
wire   [blc24ca-1:0]     hd9eac1;
wire   [blc24ca-1:0]     epab078;
wire   [blc24ca:0]       ykc1e23;
wire   [blc24ca:0]       qg788c9;
wire   [pdin_widthr-1:0]    ir23248;
wire   [pdin_widthr-1:0]    gbc9227;
wire   [pdin_widthr-1:0]    hbd80ed;
wire   [pdin_widthr-1:0]    ph3b7a;
wire   [pdin_widthr-1:0]    sue077c;
wire   [pdin_widthr-1:0]    mt1df0e;
wire   [xj71cad-1:0]    fa7c3a1;
wire   [xj71cad-1:0]    xye852;
                                                                        
            
                           ofdc411_FFTC2048            #(.by6c251(pdin_widthr),              .jp6128b(xj71cad),              .rv945f(0),              .device_family(device_family)           )         nr4a2f1 (            .clk(clk),                   .rstn(rstn),                 .ks82361(sue077c),              .hq11b09(fa7c3a1),              .mg8d84a(xw63336)                  );
      ofdc411_FFTC2048            #(.by6c251(pdin_widthr),              .jp6128b(xj71cad),              .rv945f(0),              .device_family(device_family)           )         aaa3bd9 (            .clk(clk),                   .rstn(rstn),                 .ks82361(mt1df0e),              .hq11b09(xye852),              .mg8d84a(alccd96)                  );
      ofdc411_FFTC2048            #(.by6c251(pdin_widthr),              .jp6128b(xj71cad),              .rv945f(0),              .device_family(device_family)           )         lq47d36 (            .clk(clk),                   .rstn(rstn),                 .ks82361(sue077c),              .hq11b09(xye852),              .mg8d84a(qv365ab)                  );
      ofdc411_FFTC2048            #(.by6c251(pdin_widthr),              .jp6128b(xj71cad),              .rv945f(0),              .device_family(device_family)           )         viee74e (            .clk(clk),                   .rstn(rstn),                 .ks82361(mt1df0e),              .hq11b09(fa7c3a1),              .mg8d84a(hq96aea)                  );
         generate         if(kqef411==1) begin            do9c345_FFTC2048               #(.fc2aae9(blc24ca))            ana1624               (.clk(clk), .rstn(rstn), .din(xw63336), .dout(wlaba9e));
            do9c345_FFTC2048               #(.fc2aae9(blc24ca))            qtc620c               (.clk(clk), .rstn(rstn), .din(alccd96), .dout(meea7ab));
            do9c345_FFTC2048               #(.fc2aae9(blc24ca))            mr7f2c9               (.clk(clk), .rstn(rstn), .din(qv365ab), .dout(hd9eac1));
            do9c345_FFTC2048               #(.fc2aae9(blc24ca))            vvf66bd               (.clk(clk), .rstn(rstn), .din(hq96aea), .dout(epab078));         end         else begin            assign wlaba9e = xw63336 ;            assign meea7ab = alccd96 ;            assign hd9eac1 = qv365ab ;            assign epab078 = hq96aea ;         end      endgenerate
         assign ykc1e23 = wlaba9e-meea7ab;      assign qg788c9 = hd9eac1+epab078;
         assign ir23248 = ykc1e23[gqbc4d3:kdd3134];      assign gbc9227 = qg788c9[gqbc4d3:kdd3134];
         generate         if(yx7a088==1) begin            do9c345_FFTC2048               #(.fc2aae9(pdin_widthr))            wl3979e               (.clk(clk), .rstn(rstn), .din(ir23248), .dout(hbd80ed));
            do9c345_FFTC2048               #(.fc2aae9(pdin_widthr))            qib3bf4               (.clk(clk), .rstn(rstn), .din(gbc9227), .dout(ph3b7a));
         end         else begin            assign hbd80ed = ir23248 ;            assign ph3b7a = gbc9227 ;         end      endgenerate
         generate         if(ui7de82==1) begin            do9c345_FFTC2048               #(.fc2aae9(pdin_widthr))            uk155d4               (.clk(clk), .rstn(rstn), .din(ph38443), .dout(sue077c));            do9c345_FFTC2048               #(.fc2aae9(xj71cad))            rvc956               (.clk(clk), .rstn(rstn), .din(wlbe0cb), .dout(fa7c3a1));            do9c345_FFTC2048               #(.fc2aae9(pdin_widthr))            phafd56               (.clk(clk), .rstn(rstn), .din(ri110f7), .dout(mt1df0e));            do9c345_FFTC2048               #(.fc2aae9(xj71cad))            aaa9317               (.clk(clk), .rstn(rstn), .din(zm832e8), .dout(xye852));         end         else begin            assign sue077c = ph38443 ;            assign fa7c3a1 = wlbe0cb ;            assign mt1df0e = ri110f7 ;            assign xye852 = zm832e8 ;         end      endgenerate
   endmodule                                                                                                
`timescale 1 ns / 100 ps
module sj17173_FFTC2048 (
                   clk,       
                   rstn,      
                   ibstart,   
                   points,    
                   pointset,  
                   mode,      
                   modeset,   
                   dire,      
                   diim,      
                   ibend,     
                   rfib,      
                   outvalid,  
                   obstart,   
                   except,    
                   dore,      
                   doim       
                   );
parameter pnfft_width      = 8;
parameter pdyn_points      = 0;
parameter pdin_widthr      = 16;
parameter ptwid_widthr     = 16;
parameter pdout_widthr     = 16;
parameter pnum_points      = 16;
parameter plog2_points     = 4;
parameter fixed_scaling    = 1;
parameter device_family    = "ECP";
parameter bit_reverse      = 0;
parameter rounding_method  = 1;
parameter fft_mode         = 0;
parameter pfe3535        = 0;
parameter pebr_thresh      = 7;
parameter phard_mac        = 1;
parameter pscale_reg       = 0;
parameter ptrunc_laststgs  = 0;
parameter pbfimux_level    = 0;
parameter pcntmux_level    = 0;
localparam co2b2ce      = 2*pdin_widthr;
localparam ng114ec     = 2*pdout_widthr;
localparam vve6110     = 2*ptwid_widthr;
localparam rtec748  = plog2_points-1;
localparam kf1d23b      = (plog2_points-1)/4;
localparam lq48eef      = (plog2_points-1-(4*kf1d23b))/2;
localparam fndded8          = (plog2_points-1)/2;
localparam xj7b630           = fndded8*2+1;
input                                     clk;
input                                     rstn;
input                                     ibstart;
input  [pnfft_width-1:0]                  points;
input                                     pointset;
input                                     mode;
input                                     modeset;
input  [pdin_widthr-1:0]                  dire;
input  [pdin_widthr-1:0]                  diim;
output                                    ibend;
output                                    rfib;
output                                    outvalid;
output                                    obstart;
output                                    except;
output [pdout_widthr-1:0]                 dore;
output [pdout_widthr-1:0]                 doim;
wire                                      clk;
wire                                      rstn;
wire                                      ibstart;
wire                                      outvalid;
wire                                      obstart;
wire  [pdin_widthr-1:0]                   dire;
wire  [pdin_widthr-1:0]                   diim;
wire                                      kq439ac;
wire                                      cm599c8;
wire                                      jc52b77;
wire  [pdin_widthr-1:0]                   kd44c3b;
wire  [pdin_widthr-1:0]                   do30eec;
wire  [pdin_widthr-1:0]                   ec3bb19;
wire  [pdin_widthr-1:0]                   zxec646;
wire                                      ir95bbb;
wire  [pdout_widthr-1:0]                  ldc8dd7;
wire  [pdout_widthr-1:0]                  rv375f8;
wire  [pdout_widthr-1:0]                  pfd7e3e;
wire  [pdout_widthr-1:0]                  wjf8fbf;
wire                                      ribd9a1;
wire                                      ho5224c;
wire                                      ph91262;
wire                                      do89317;
wire  [pdin_widthr-1:0]                   cm498ba;
wire  [pdin_widthr-1:0]                   yk4c5d1;
wire  [pnfft_width-1:0]                   ksbc8fe;
wire  [plog2_points:0]                    an39028;
wire  [plog2_points:0]                    pfcdf4c;
wire  [plog2_points-1:0]                  mt12817;
wire  [plog2_points:0]                    qgeff2b;
wire  [plog2_points:0]                    fnc8144;
wire  [plog2_points:0]                    kdf8b37;
wire  [plog2_points+1:0]                  je2a081;
wire  [plog2_points+1:0]                  os67205;
wire  [plog2_points*(plog2_points+1)-1:0] bn289b8;
wire  [co2b2ce*(plog2_points+2)-1:0]  ofc9c10;
wire  [vve6110*(plog2_points+1)-1:0] wwe5667;
wire  [pdout_widthr*2-1:0]                tw35837;
wire  [co2b2ce-1:0]                   yx7f959;
wire                                      vkb84a0;
wire                                      rtc2502;
wire                                      lsbdfe5;
wire  [plog2_points:0]                    qi5137;
wire                                      wla1295;
wire                                      of54252;
wire                                      ymac1bb;
wire     os78568;
wire     ou2b339;
genvar rtd7680,qvbb406,hq869c2,pf40c19;
wire[`TWID_WIDTH-1:0]   dme1d4e;
wire[`TWID_WIDTH-1:0]   wj75392;
                                                                                                                  
                                                   assign os78568 = rfib & ibstart ;
                     uifa97e_FFTC2048 osfa795 (            .clk            (clk),                        .rstn           (rstn),                                   .ibstart        (os78568),                    .modeset        (modeset),                    .mode           (mode),           
            .wl80cf8          (jc52b77)                   );
         generate      begin         if (pdyn_points==1) begin         db947c_FFTC2048 #(                    .plog2_points(plog2_points),                    .pbfimux_level     (pbfimux_level),                    .pcntmux_level     (pcntmux_level),                    .pnfft_width(pnfft_width))            vk4cf4 (            .clk      (clk),                   .rstn     (rstn),                  .ibstart  (os78568),               .points   (points),                .pointset (pointset),              .kdf8b37      ({(plog2_points+1){1'b0}}),            .ksbc8fe  (ksbc8fe),               .mt12817    (mt12817),                 .lsbdfe5(lsbdfe5),             .wla1295(wla1295),            .sw1fc5d(),            .jcc59bd     (),            .qgeff2b   (qgeff2b)     
            );         end         else begin            assign  ksbc8fe   = 0;            assign  mt12817     = 0;            assign  lsbdfe5 = 1'b0;            assign  qgeff2b    = 0;            assign  wla1295= 1'b0;         end      end      endgenerate
         defparam kq6d7ae.fc2aae9=pdin_widthr;
      gdd98d_FFTC2048 kq6d7ae (            .clk            (clk),                        .rstn           (rstn),                       .ibstart        (os78568),                    .dire           (dire),                       .diim           (diim),                       .ribd9a1       (ribd9a1),                   .ho5224c      (ho5224c),                  .ph91262      (ph91262),                  .do89317      (do89317),                  .cm498ba          (cm498ba),                      .yk4c5d1          (yk4c5d1)                       );
            assign kd44c3b = cm498ba;         assign do30eec = yk4c5d1;
         aabcb24_FFTC2048         #(                     .fc2aae9(pdin_widthr),                     .ls89b60(0))              uv605dc (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .fft_mode      (jc52b77     ),                     .ec24226        (              ),                     .dire          (kd44c3b      ),                     .diim          (do30eec      ),                     .dore          (ec3bb19      ),                     .doim          (zxec646      )                 );
      assign ofc9c10[co2b2ce-1:0]    = {ec3bb19,zxec646};      assign je2a081[0]                  = 1'b0;      assign rtc2502                 =je2a081[0];      assign yx7f959                  = {ec3bb19,zxec646};
      generate      begin         if (pscale_reg==1) begin            assign kdf8b37[0]            = ph91262;            assign vkb84a0           = do89317;                                 end         else begin            assign kdf8b37[0]            = ho5224c;            assign vkb84a0           = ph91262;         end      end      endgenerate
         generate      begin         for (rtd7680=0; rtd7680<plog2_points; rtd7680=rtd7680+1) begin:vvfc975            ls1e5c2_FFTC2048  #(                  .pdyn_points       (pdyn_points),                  .plog2_points(plog2_points),                  .twb8d6f(rtd7680),                  .enc6b7b(pdin_widthr),                  .hq35bdc(plog2_points-(rtd7680+1)),                  .hqadee3(fixed_scaling),                  .rounding_method   (rounding_method),                  .ptwid_widthr(ptwid_widthr),                  .pfe3535(pfe3535),                  .xj7b8d4(plog2_points),                  .gq1a9ae((plog2_points-rtd7680-1)/pebr_thresh),                  .med4d71(device_family),                  .pscale_reg(pscale_reg),                  .ptrunc_laststgs   (ptrunc_laststgs),                  .vv7105c      (bit_reverse),                  .phard_mac(phard_mac)                  )                the3a30 (                  .clk           (clk),                                                             .rstn          (rstn),                                                            .vkb84a0       (vkb84a0),                                                         .rtc2502       (rtc2502),                                                         .mt12817         (mt12817),                                                           .lsbdfe5     (lsbdfe5),                                                       .hd940bd        (kdf8b37[rtd7680]),                                                          .tja05ef        (kdf8b37[rtd7680+1]),                                                        .sj2f7f        (je2a081[rtd7680]),                                                          .qv17bfc        (je2a081[rtd7680+1]),                                                        .ou2b339      (ou2b339),                                                        .cm599c8      (cm599c8),                                                        .encce40     (os67205[rtd7680+1]),                                                   .os67205      (os67205[rtd7680]),                                                     .fnc8144          (fnc8144[rtd7680+1]),                                                       .an39028  (an39028[rtd7680+1]),                                               .vv40a26     (pfcdf4c[rtd7680+1]),                                                    .qi5137           (qi5137[rtd7680+1]),                                                       .qgeff2b        (qgeff2b[rtd7680]),                                                       .yx7f959        (yx7f959),                                                          .pffcacc           (ofc9c10[co2b2ce*(rtd7680+1)-1:co2b2ce*rtd7680]),                          .bn289b8         (bn289b8[plog2_points*(rtd7680+2)-1:plog2_points*(rtd7680+1)]),                  .wwe5667           (wwe5667[vve6110*(rtd7680+2)-1:vve6110*(rtd7680+1)]),                    .en44dc6          (ofc9c10[co2b2ce*(rtd7680+2)-1:co2b2ce*(rtd7680+1)])                       );         end      end      endgenerate   
         
      generate      begin         for(qvbb406=2;qvbb406<plog2_points;qvbb406=qvbb406+2) begin:kde26ef            if(qvbb406==2) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid0FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==4) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid1FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==6) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid2FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==8) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid3FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==10) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid4FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==12) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid5FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==14) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid6FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end         end      end      endgenerate
   
         defparam eac1326.bit_reverse    = bit_reverse;      defparam eac1326.plog2_points   = plog2_points;      defparam eac1326.enc6b7b   = pdout_widthr;      defparam eac1326.pdyn_points    = pdyn_points;      defparam eac1326.pnfft_width    = pnfft_width;      defparam eac1326.med4d71 = device_family;
      ale81d9_FFTC2048 eac1326 (            .clk                (clk),                                                                        .rstn               (rstn),                                                                       .qi5137                (qi5137),                                                                        .an39028       (an39028),                                                               .pfcdf4c          (pfcdf4c),                                                                  .os67205           (os67205),                                                                  .mt12817              (mt12817),                                                                      .lsbdfe5          (lsbdfe5),                                                                  .kq4cf46             (fnc8144[plog2_points-1]),                                                       .kq67a31           (kdf8b37[plog2_points-1]),                                                        .zz3d189            (ofc9c10[co2b2ce*(plog2_points)-1:co2b2ce*(plog2_points-1)]),             .fnc8144               (fnc8144[plog2_points]),                                                                     .ip75347                (of54252),            .hd940bd             (kdf8b37[plog2_points]),                                                          .ri89d08              (ofc9c10[co2b2ce*(plog2_points+1)-1:co2b2ce*plog2_points]),               .ksbc8fe            (ksbc8fe),                                                                    .except             (except),                                                                     .ou2b339           (ou2b339),                                                                   .outvalid           (outvalid),                                                                   .kq439ac           (kq439ac),                                                                   .cm599c8           (cm599c8),                                                                   .obstart            (obstart),                                                                    .tw35837             (tw35837),                                                                     .ymac1bb         (ymac1bb)            );
            assign ldc8dd7 = tw35837[pdout_widthr*2-1:pdout_widthr];         assign rv375f8 = tw35837[pdout_widthr-1:0];
         aabcb24_FFTC2048         #(                     .fc2aae9(pdout_widthr),                     .ls89b60(1))              oh17611 (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .fft_mode      (ir95bbb     ),                     .ec24226        (ymac1bb    ),                     .dire          (ldc8dd7      ),                     .diim          (rv375f8      ),                     .dore          (pfd7e3e      ),                     .doim          (wjf8fbf      )                 );
         assign dore = pfd7e3e;      assign doim = wjf8fbf;            
         defparam qi97f50.bit_reverse=bit_reverse;      defparam qi97f50.pdyn_points=pdyn_points;      wwdbe0f_FFTC2048 qi97f50 (            .clk            (clk),                        .rstn           (rstn),                       .mec1e54       (os78568),                    .ibstart        (ribd9a1),                   .os67205       (os67205[0]),                .qi5137            (qi5137[plog2_points]),            .of54252        (of54252),            .wla1295     (wla1295),            .rv94ad (kdf8b37[plog2_points]),            .cm599c8       (kq439ac),                   .jc52b77      (jc52b77     ),            .ir95bbb      (ir95bbb     ),            .ibend          (ibend),                      .rfib           (rfib)                        );
   endmodule                                                                                                
`timescale 1 ns / 100 ps
module al4458b_FFTC2048 (
                   clk,       
                   rstn,      
                   ibstart,   
                   points,    
                   pointset,  
                   mode,      
                   modeset,   
                   sfact,     
                   sfactset,  
                   dire,      
                   diim,      
                   ibend,     
                   rfib,      
                   outvalid,  
                   obstart,   
                   except,    
                   dore,      
                   doim       
                   );
parameter pnfft_width      = 8;
parameter pdyn_points      = 0;
parameter pdin_widthr      = 16;
parameter ptwid_widthr     = 16;
parameter pdout_widthr     = 16;
parameter pnum_points      = 16;
parameter plog2_points     = 4;
parameter fixed_scaling    = 1;
parameter device_family    = "ECP";
parameter bit_reverse      = 0;
parameter sfact_width      = 16;
parameter rounding_method  = 1;
parameter fft_mode         = 0;
parameter pfe3535        = 0;
parameter pebr_thresh      = 7;
parameter phard_mac        = 1;
parameter pscale_reg       = 0;
parameter ptrunc_laststgs  = 0;
parameter pbfimux_level    = 0;
parameter pcntmux_level    = 0;
localparam co2b2ce      = 2*pdin_widthr;
localparam ng114ec     = 2*pdout_widthr;
localparam vve6110     = 2*ptwid_widthr;
localparam rtec748  = plog2_points-1;
localparam kf1d23b      = (plog2_points-1)/4;
localparam lq48eef      = (plog2_points-1-(4*kf1d23b))/2;
localparam fndded8          = (plog2_points-1)/2;
localparam xj7b630           = fndded8*2+1;
input                                     clk;
input                                     rstn;
input                                     ibstart;
input  [pnfft_width-1:0]                  points;
input                                     pointset;
input                                     mode;
input                                     modeset;
input  [sfact_width-1:0]                  sfact;
input                                     sfactset;
input  [pdin_widthr-1:0]                  dire;
input  [pdin_widthr-1:0]                  diim;
output                                    except;
output                                    ibend;
output                                    rfib;
output                                    outvalid;
output                                    obstart;
output [pdout_widthr-1:0]                 dore;
output [pdout_widthr-1:0]                 doim;
wire                                      clk;
wire                                      rstn;
wire                                      ibstart;
wire                                      outvalid;
wire                                      obstart;
wire  [pdin_widthr-1:0]                   dire;
wire  [pdin_widthr-1:0]                   diim;
wire                                      kq439ac;
wire                                      cm599c8;
wire                                      jc52b77;
wire  [pdin_widthr-1:0]                   kd44c3b;
wire  [pdin_widthr-1:0]                   do30eec;
wire  [pdin_widthr-1:0]                   ec3bb19;
wire  [pdin_widthr-1:0]                   zxec646;
wire                                      ir95bbb;
wire  [pdout_widthr-1:0]                  ldc8dd7;
wire  [pdout_widthr-1:0]                  rv375f8;
wire  [pdout_widthr-1:0]                  pfd7e3e;
wire  [pdout_widthr-1:0]                  wjf8fbf;
wire                                      ph91262;
wire                                      ho5224c;
wire                                      do89317;
wire                                      ribd9a1;
wire  [pdin_widthr-1:0]                   cm498ba;
wire  [pdin_widthr-1:0]                   yk4c5d1;
wire  [pnfft_width-1:0]                   ksbc8fe;
wire  [plog2_points:0]                    an39028;
wire  [plog2_points:0]                    pfcdf4c;
wire  [plog2_points-1:0]                  mt12817;
wire  [plog2_points:0]                    qgeff2b;
wire  [plog2_points:0]                    fnc8144;
wire  [plog2_points:0]                    kdf8b37;
wire  [plog2_points:0]                    sw1fc5d;
wire  [plog2_points+1:0]                  je2a081;
wire  [plog2_points+1:0]                  os67205;
wire  [plog2_points*(plog2_points+1)-1:0] bn289b8;
wire  [vve6110*(plog2_points+1)-1:0] wwe5667;
wire  [(plog2_points+2)*(plog2_points+1)+co2b2ce*(plog2_points+2)-1:0]  ofc9c10;
wire  [pdout_widthr*2-1:0]                tw35837;
wire  [sfact_width-1:0]                   an2cdeb;
wire  [co2b2ce-1:0]                   sh414c9;
wire  [ng114ec-1:0]                  yx7f959;
wire                                      vkb84a0;
wire                                      rtc2502;
wire                                      lsbdfe5;
wire  [pdout_widthr-1:0]                  yz8747;
wire  [pdout_widthr-1:0]                  kf1d1e0;
wire  [pdin_widthr-1+plog2_points:0]      ux3c162;
wire  [pdin_widthr-1+plog2_points:0]      yz2c501;
wire                                      jcc59bd;
wire  [plog2_points:0]                    qi5137;
wire                                      wla1295;
wire                                      of54252;
wire                                      ymac1bb;
wire     os78568;
wire                                      ou2b339;
genvar rtd7680,qvbb406,hq869c2,pf40c19;
wire[`TWID_WIDTH-1:0]   dme1d4e;
wire[`TWID_WIDTH-1:0]   wj75392;
                                                                                                                        
                                                   assign os78568 = rfib & ibstart ;
            
         uifa97e_FFTC2048 osfa795 (            .clk            (clk),                        .rstn           (rstn),                                   .ibstart        (os78568),                    .modeset        (modeset),                    .mode           (mode),           
            .wl80cf8          (jc52b77)                   );
         defparam gd2cb1.sfact_width=sfact_width;      defparam gd2cb1.plog2_points = plog2_points;      defparam gd2cb1.pdyn_points = pdyn_points;
      ph1c7c6_FFTC2048 gd2cb1 (            .clk            (clk),                        .rstn           (rstn),                                   .ibstart        (os78568),                    .sfact          (sfact),                      .sfactset       (sfactset),                   .kdf8b37            (sw1fc5d),            .jcc59bd           (jcc59bd),                        .lsbdfe5(lsbdfe5), 
            .an2cdeb         (an2cdeb)                      );
         generate      begin         if (pdyn_points==1) begin         db947c_FFTC2048 #(                    .plog2_points(plog2_points),                    .pbfimux_level     (pbfimux_level),                    .pcntmux_level     (pcntmux_level),                    .pnfft_width(pnfft_width))            vk4cf4 (            .clk      (clk),                   .rstn     (rstn),                  .ibstart  (os78568),               .points   (points),                .pointset (pointset),              .kdf8b37      (kdf8b37),            .ksbc8fe  (ksbc8fe),               .mt12817    (mt12817),                 .lsbdfe5(lsbdfe5),             .wla1295(wla1295),            .sw1fc5d(sw1fc5d),            .jcc59bd     (jcc59bd),            .qgeff2b   (qgeff2b)     
            );         end         else begin            assign  ksbc8fe   = 0;            assign  mt12817     = 0;            assign  lsbdfe5 = 1'b0;            assign  qgeff2b    = 0;            assign  sw1fc5d = kdf8b37;            assign  jcc59bd      = kdf8b37[1];            assign  wla1295= 1'b0;         end      end      endgenerate
         defparam kq6d7ae.fc2aae9=pdin_widthr;
      gdd98d_FFTC2048 kq6d7ae (            .clk            (clk),                        .rstn           (rstn),                       .ibstart        (os78568),                    .dire           (dire),                       .diim           (diim),                       .ribd9a1       (ribd9a1),                   .ho5224c      (ho5224c),                  .ph91262      (ph91262),                  .do89317      (do89317),                  .cm498ba          (cm498ba),                      .yk4c5d1          (yk4c5d1)                       );            
            assign kd44c3b = cm498ba;         assign do30eec = yk4c5d1;
         aabcb24_FFTC2048         #(                     .fc2aae9(pdin_widthr),                     .ls89b60(0))              uv605dc (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .fft_mode      (jc52b77     ),                     .ec24226        (              ),                     .dire          (kd44c3b      ),                     .diim          (do30eec      ),                     .dore          (ec3bb19      ),                     .doim          (zxec646      )                 );                 
      assign ofc9c10[co2b2ce-1:0]    = {ec3bb19,zxec646};      assign je2a081[0]                  = 1'b0;      assign rtc2502                 =je2a081[0];
      assign yz2c501                 ={{plog2_points{zxec646[pdin_widthr-1]}},zxec646};      assign ux3c162                 ={{plog2_points{ec3bb19[pdin_widthr-1]}},ec3bb19};
      generate      begin         if (pscale_reg==1) begin            assign kdf8b37[0]            = ph91262;            assign vkb84a0           = do89317;                                 end         else begin            assign kdf8b37[0]            = ho5224c;            assign vkb84a0           = ph91262;         end      end      endgenerate
         generate      begin         for (rtd7680=0; rtd7680<plog2_points; rtd7680=rtd7680+1) begin:vvfc975                        me68523_FFTC2048  #(                  .pdyn_points       (pdyn_points),                  .plog2_points(plog2_points),                  .twb8d6f(rtd7680),                  .enc6b7b(pdin_widthr+rtd7680),                  .hq35bdc(plog2_points-(rtd7680+1)),                  .hqadee3(fixed_scaling),                  .rounding_method   (rounding_method),                  .ptwid_widthr(ptwid_widthr),                  .pfe3535(pfe3535),                  .xj7b8d4(plog2_points),                  .gq1a9ae((plog2_points-rtd7680-1)/pebr_thresh),                  .med4d71(device_family),                  .phard_mac(phard_mac),                  .pscale_reg(pscale_reg),                  .ptrunc_laststgs   (ptrunc_laststgs),                  .vv7105c      (bit_reverse),                  .xyadfc4(pdin_widthr)                  )                the3a30 (                  .clk           (clk),                  .rstn          (rstn),                  .vkb84a0       (vkb84a0),                                                         .rtc2502       (rtc2502),                                                         .mt12817         (mt12817),                                                           .lsbdfe5     (lsbdfe5),                                                       .hd940bd        (kdf8b37[rtd7680]),                  .tja05ef        (kdf8b37[rtd7680+1]),                  .sj2f7f        (je2a081[rtd7680]),                  .aaacedc        (an2cdeb[2*plog2_points-1-(2*rtd7680+0):2*plog2_points-1-(2*rtd7680+1)]),                  .qv17bfc        (je2a081[rtd7680+1]),                  .ou2b339      (ou2b339),                                                        .cm599c8      (cm599c8),                                                        .encce40     (os67205[rtd7680+1]),                                                   .os67205      (os67205[rtd7680]),                  .fnc8144          (fnc8144[rtd7680+1]),                  .an39028  (an39028[rtd7680+1]),                                               .vv40a26     (pfcdf4c[rtd7680+1]),                                                    .qi5137           (qi5137[rtd7680+1]),                                                       .qgeff2b        (qgeff2b[rtd7680]),                                                                                                             .yx7f959        ({ux3c162[pdin_widthr+rtd7680-1:0],yz2c501[pdin_widthr+rtd7680-1:0]}),                   .pffcacc           (ofc9c10[(rtd7680+1)*rtd7680+co2b2ce*(rtd7680+1)-1:rtd7680*(rtd7680-1)+co2b2ce*rtd7680]),                  .bn289b8         (bn289b8[plog2_points*(rtd7680+2)-1:plog2_points*(rtd7680+1)]),                  .wwe5667           (wwe5667[vve6110*(rtd7680+2)-1:vve6110*(rtd7680+1)]),                  .en44dc6          (ofc9c10[(rtd7680+2)*(rtd7680+1)+co2b2ce*(rtd7680+2)-1:(rtd7680+1)*rtd7680+co2b2ce*(rtd7680+1)])                  );         end      end      endgenerate
      generate      begin         for(qvbb406=2;qvbb406<plog2_points;qvbb406=qvbb406+2) begin:kde26ef            if(qvbb406==2) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid0FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==4) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid1FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==6) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid2FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==8) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid3FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==10) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid4FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==12) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid5FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end else if(qvbb406==14) begin               tue1eff_FFTC2048 #(                        .qgfa399      (plog2_points-qvbb406+2  ),                        .ead1cc9      (`TWID_WIDTH   ),                        .rv8e648     ("reg"       ),                        .ps73247   ("twid6FFTC2048.mem"    ),                        .tw9923b      (device_family ),                        .ofc91db        (2             ),                        .ne48edc       (1024          ))               suf55ba (                        .rstn    (rstn    ),                        .clk     (clk     ),                        .bydfe8e   (bn289b8[plog2_points*(qvbb406+2)-1:plog2_points*(qvbb406+1)+(qvbb406-2)]),                        .dout    (wwe5667[vve6110*(qvbb406+2)-1:vve6110*(qvbb406+1)])                     );            end         end      end      endgenerate
   
      assign   kf1d1e0 = {ofc9c10[pdout_widthr-2+(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1)],ofc9c10[pdout_widthr-2+(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1):(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1)]};      assign   yz8747 = {ofc9c10[pdout_widthr*2-3+(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1)],ofc9c10[pdout_widthr*2-3+(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1):pdout_widthr-1+(plog2_points-1)*(plog2_points-2)+co2b2ce*(plog2_points-1)]};
         defparam eac1326.bit_reverse    = bit_reverse;      defparam eac1326.plog2_points   = plog2_points;      defparam eac1326.enc6b7b   = pdout_widthr;      defparam eac1326.pdyn_points    = pdyn_points;      defparam eac1326.pnfft_width    = pnfft_width;      defparam eac1326.med4d71 = device_family;
      ale81d9_FFTC2048 eac1326 (            .clk      (clk),            .rstn     (rstn),            .qi5137                (qi5137),                                                    .an39028       (an39028),                                           .pfcdf4c          (pfcdf4c),                                              .os67205           (os67205),                                               .mt12817              (mt12817),                                                  .lsbdfe5          (lsbdfe5),                                              .kq4cf46             (fnc8144[plog2_points-1]),                                   .kq67a31           (kdf8b37[plog2_points-1]),                                                            .zz3d189            ({yz8747,kf1d1e0}),                                  .fnc8144     (fnc8144[plog2_points]),                        .ip75347      (of54252),            .hd940bd   (kdf8b37[plog2_points]),            .ri89d08    (ofc9c10[(plog2_points+1)*plog2_points+co2b2ce*(plog2_points+1)-1:plog2_points*(plog2_points-1)+co2b2ce*plog2_points]),            .ksbc8fe  (ksbc8fe),                                                          .except   (except),                                                           .ou2b339 (ou2b339),                                                         .outvalid (outvalid),            .kq439ac (kq439ac),            .cm599c8 (cm599c8),                                                         .obstart  (obstart),            .tw35837   (tw35837),            .ymac1bb(ymac1bb)            );
         assign ldc8dd7 = tw35837[pdout_widthr*2-1:pdout_widthr];      assign rv375f8 = tw35837[pdout_widthr-1:0];
      aabcb24_FFTC2048 #(            .fc2aae9(pdout_widthr),            .ls89b60(1))         oh17611 (            .clk           (clk           ),            .rstn          (rstn          ),            .fft_mode      (ir95bbb     ),            .ec24226        (ymac1bb    ),            .dire          (ldc8dd7      ),            .diim          (rv375f8      ),            .dore          (pfd7e3e      ),            .doim          (wjf8fbf      )            );
         assign dore = pfd7e3e;      assign doim = wjf8fbf;            
         defparam qi97f50.bit_reverse=bit_reverse;      defparam qi97f50.pdyn_points=pdyn_points;      wwdbe0f_FFTC2048 qi97f50 (            .clk            (clk),                        .rstn           (rstn),                       .mec1e54       (os78568),                    .ibstart        (ribd9a1),                      .os67205       (os67205[0]),                .qi5137            (qi5137[plog2_points]),            .of54252        (of54252),                      .wla1295     (wla1295),                   .rv94ad (kdf8b37[plog2_points]),            .cm599c8       (kq439ac),                   .jc52b77      (jc52b77     ),             .ir95bbb      (ir95bbb     ),             .ibend          (ibend),                      .rfib           (rfib)                        );
   endmodule                                                                                                
`timescale 1 ns / 100 ps
module twbd919_FFTC2048 (
                   clk,       
                   rstn,      
                   ibstart,   
                   points,    
                   pointset,  
                   mode,      
                   modeset,   
                   sfact,     
                   sfactset,  
   
                   dire,      
                   diim,      
                   ibend,     
                   rfib,      
                   outvalid,  
                   obstart,   
                   except,    
                   dore,      
                   doim       
                   );
parameter pnfft_width      = 8;
parameter pdyn_points      = 0;
parameter pdin_widthr      = 16;
parameter ptwid_widthr     = 16;
parameter pdout_widthr     = 16;
parameter pnum_points      = 16;
parameter plog2_points     = 4;
parameter fixed_scaling    = 1;
parameter device_family    = "ECP";
parameter bit_reverse      = 0;
parameter sfact_width      = 16;
parameter rounding_method  = 1;
parameter fft_mode         = 0;
parameter pfe3535        = 0;
parameter pebr_thresh      = 7;
parameter phard_mac        = 1;
parameter pscale_reg       = 0;
parameter ptrunc_laststgs  = 0;
parameter pbfimux_level    = 0;
parameter pcntmux_level    = 0;
input                                     clk;
input                                     rstn;
input                                     ibstart;
input  [pnfft_width-1:0]                  points;
input                                     pointset;
input                                     mode;
input                                     modeset;
input  [sfact_width-1:0]                  sfact;
input                                     sfactset;
input  [pdin_widthr-1:0]                  dire;
input  [pdin_widthr-1:0]                  diim;
output                                    ibend;
output                                    rfib;
output                                    outvalid;
output                                    obstart;
output                                    except;
output [pdout_widthr-1:0]                 dore;
output [pdout_widthr-1:0]                 doim;
wire                                      clk;
wire                                      rstn;
wire                                      ibstart;
wire                                      outvalid;
wire                                      obstart;
wire  [pdin_widthr-1:0]                   dire;
wire  [pdin_widthr-1:0]                   diim;
wire                                      ribd9a1;
wire  [pdin_widthr-1:0]                   cm498ba;
wire  [pdin_widthr-1:0]                   yk4c5d1;
                                                                                                                        
                           
   generate      if (( fixed_scaling==0 ) || ( fixed_scaling==3 )) begin          al4458b_FFTC2048 #(            .pnfft_width       (pnfft_width),            .pdyn_points       (pdyn_points),            .pdin_widthr       (pdin_widthr),            .ptwid_widthr      (ptwid_widthr),            .pdout_widthr      (pdout_widthr),            .pnum_points       (pnum_points),            .plog2_points      (plog2_points),            .fixed_scaling     (fixed_scaling),            .rounding_method   (rounding_method),            .device_family     (device_family),            .bit_reverse       (bit_reverse),            .fft_mode          (fft_mode),            .pfe3535         (pfe3535),            .sfact_width       (sfact_width),            .pebr_thresh       (pebr_thresh),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .pbfimux_level     (pbfimux_level),            .pcntmux_level     (pcntmux_level),            .phard_mac         (phard_mac)            )           nt27f5f (            .clk               (clk),                     .rstn              (rstn),                    .ibstart           (ibstart),                 .pointset          (pointset),                .points            (points),                  .modeset           (modeset),                 .mode              (mode),                    .sfact             (sfact),                   .sfactset          (sfactset),                .dire              (dire),                    .diim              (diim),                    .ibend             (ibend),                   .rfib              (rfib),                    .outvalid          (outvalid),                .obstart           (obstart),                 .except            (except),                  .dore              (dore),                    .doim              (doim)                     );      end      else begin         sj17173_FFTC2048 #(            .pnfft_width       (pnfft_width),            .pdyn_points       (pdyn_points),            .pdin_widthr       (pdin_widthr),            .ptwid_widthr      (ptwid_widthr),            .pdout_widthr      (pdout_widthr),            .pnum_points       (pnum_points),            .plog2_points      (plog2_points),            .fixed_scaling     (fixed_scaling),            .rounding_method   (rounding_method),            .bit_reverse       (bit_reverse),            .fft_mode          (fft_mode),            .pfe3535         (pfe3535),            .device_family     (device_family),            .pebr_thresh       (pebr_thresh),            .pscale_reg        (pscale_reg),            .ptrunc_laststgs   (ptrunc_laststgs),            .pbfimux_level     (pbfimux_level),            .pcntmux_level     (pcntmux_level),            .phard_mac         (phard_mac)            )           ne4d871 (            .clk               (clk),                     .rstn              (rstn),                    .ibstart           (ibstart),                 .pointset          (pointset),                .points            (points),                  .modeset           (modeset),                 .mode              (mode),                    .dire              (dire),                    .diim              (diim),                    .ibend             (ibend),                   .rfib              (rfib),                    .outvalid          (outvalid),                .obstart           (obstart),                 .except            (except),                  .dore              (dore),                    .doim              (doim)                     );      end   endgenerate
   endmodule
`else
                                                                                          
`timescale 1 ns / 100 ps
module rt550ab_FFTC2048(
             clk,                       
             rstn,                      
             mg157da,                
             gdabed1,                
             xj5f68d,                
             psfb46e,                
             xwda373,               
             osd1b9a,               
             qi8dcd0,               
             jp6e681                
            ) ;
parameter   ps7340e = 8;
input                      clk ;
input                      rstn ;
input [ps7340e-1:0]     mg157da ;
input [ps7340e-1:0]     gdabed1 ;
input [ps7340e-1:0]     xj5f68d ;
input [ps7340e-1:0]     psfb46e ;
output[ps7340e:0]       xwda373 ;
output[ps7340e:0]       osd1b9a ;
output[ps7340e:0]       qi8dcd0 ;
output[ps7340e:0]       jp6e681 ;
wire[ps7340e:0]         ux29433;
wire[ps7340e:0]         zx50cef;
wire[ps7340e:0]         oh33bf3;
wire[ps7340e:0]         icefce0;
            assign ux29433 = {mg157da[ps7340e-1],mg157da};      assign zx50cef = {xj5f68d[ps7340e-1],xj5f68d};      assign oh33bf3 = {gdabed1[ps7340e-1],gdabed1};      assign icefce0 = {psfb46e[ps7340e-1],psfb46e};
            su566ea_FFTC2048 #(.wyb3750    ("ADD"            ),                  .ps7340e (ps7340e+1     ),                  .ayea07f (`DEVICE_FAMILY),                  .xj503f8  (`ADDER_PIPELINE+1))      rv81fc7 (               .rstn    (rstn          ),               .clk     (clk           ),               .ba3f16e       (ux29433       ),               .fac5b9d       (oh33bf3       ),               .jp6e75e       (xwda373   )            );
            su566ea_FFTC2048 #(.wyb3750    ("ADD"            ),                  .ps7340e (ps7340e+1     ),                  .ayea07f (`DEVICE_FAMILY),                  .xj503f8  (`ADDER_PIPELINE+1))      jr8bbdf (               .rstn    (rstn          ),               .clk     (clk           ),               .ba3f16e       (zx50cef       ),               .fac5b9d       (icefce0       ),               .jp6e75e       (qi8dcd0   )            );
            su566ea_FFTC2048 #(.wyb3750    ("SUB"            ),                  .ps7340e (ps7340e+1     ),                  .ayea07f (`DEVICE_FAMILY),                  .xj503f8  (`ADDER_PIPELINE+1))      kdf770e (               .rstn    (rstn          ),               .clk     (clk           ),               .ba3f16e       (ux29433       ),               .fac5b9d       (oh33bf3       ),               .jp6e75e       (osd1b9a   )            );
            su566ea_FFTC2048 #(.wyb3750    ("SUB"            ),                  .ps7340e (ps7340e+1     ),                  .ayea07f (`DEVICE_FAMILY),                  .xj503f8  (`ADDER_PIPELINE+1))      ea56449 (               .rstn    (rstn          ),               .clk     (clk           ),               .ba3f16e       (zx50cef       ),               .fac5b9d       (icefce0       ),               .jp6e75e       (jp6e681   )            );
   endmodule                                                                                          
`timescale 1 ns / 100 ps
module ec10059_FFTC2048(
             clk,                   
             rstn,                  
             pub262,            
             yk59313,            
             czc9899,            
             yk4c4cd,            
             os62668,            
             bn13340,            
             ri99a06,           
             vvcd032,           
             qg68196,           
             zx40cb1            
            ) ;
parameter zz658f = `BE_PL_DEPTH;
input                      clk ;
input                      rstn ;
input [`DATA_WIDTH-1:0]    pub262 ;
input [`DATA_WIDTH-1:0]    yk59313 ;
input [`DATA_WIDTH-1:0]    czc9899 ;
input [`DATA_WIDTH-1:0]    yk4c4cd ;
input [`TWID_WIDTH-1:0]    os62668 ;
input [`TWID_WIDTH-1:0]    bn13340 ;
output[`DATA_WIDTH+1:0]    ri99a06 ;
output[`DATA_WIDTH+1:0]    vvcd032 ;
output[`DATA_WIDTH+1:0]    qg68196 ;
output[`DATA_WIDTH+1:0]    zx40cb1 ;
wire[`DATA_WIDTH:0]        pse41ee ;
wire[`DATA_WIDTH:0]        ls20f73 ;
wire[`DATA_WIDTH:0]        cb7b9a ;
wire[`DATA_WIDTH:0]        tj3dcd4 ;
      dmee6a7_FFTC2048  tu7353a (                  .clk  (clk           ),                  .rstn (rstn          ),                  .ba3f16e    (yk59313    ),                  .fac5b9d    (os62668    ),                  .jp6e75e    (yk4c4cd    ),                  .pfe9af9    (bn13340    ),                  .rt6be72    (ls20f73  )                  ) ;
      thf9cbe_FFTC2048  cmce5f7 (                  .clk  (clk           ),                  .rstn (rstn          ),                  .ba3f16e    (yk59313    ),                  .fac5b9d    (bn13340    ),                  .jp6e75e    (yk4c4cd    ),                  .pfe9af9    (os62668    ),                  .rt6be72    (tj3dcd4)                  ) ;
      lqee0f9_FFTC2048 #(.gb707ca  (zz658f     ),                  .mg1f2a2 (`DATA_WIDTH+1)               ) hbf9510(                  .clk  (clk                                      ),                  .rstn (rstn                                     ),                  .pfe9af9    ({pub262[`DATA_WIDTH-1], pub262}  ),                  .hdaa0f5    (pse41ee                             )               ) ;
      lqee0f9_FFTC2048 #(.gb707ca  (zz658f     ),                  .mg1f2a2 (`DATA_WIDTH+1)               ) os774cd(                  .clk  (clk                                      ),                  .rstn (rstn                                     ),                  .pfe9af9    ({czc9899[`DATA_WIDTH-1], czc9899}  ),                  .hdaa0f5    (cb7b9a                             )               ) ;
            rt550ab_FFTC2048 #(`DATA_WIDTH+1) xy96572(                .clk          (clk           ),                .rstn         (rstn          ),                .mg157da   (pse41ee  ),                .xj5f68d   (cb7b9a  ),                .gdabed1   (ls20f73  ),                .psfb46e   (tj3dcd4  ),                .xwda373  (ri99a06   ),                .osd1b9a  (vvcd032   ),                .qi8dcd0  (qg68196   ),                .jp6e681  (zx40cb1   )               ) ;
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module su566ea_FFTC2048( rstn,
                     clk,
                     ba3f16e,
                     fac5b9d,
                     jp6e75e
                  );
parameter   wyb3750 = "ADD";
parameter   ps7340e = 8;
parameter   xj503f8 = 1;
parameter   ayea07f="ECP2";
parameter ks348d2 = ps7340e/2;
parameter sj2348d = ps7340e/2+(ps7340e%2);
input                   rstn;
input                   clk;
input [ps7340e-1:0]  ba3f16e;
input [ps7340e-1:0]  fac5b9d;
output[ps7340e-1:0]  jp6e75e;
wire[ps7340e-1:0] pfe6b30;
wire[sj2348d-1:0]  mgacc3b;
wire[sj2348d-1:0]  ri30ec2;
wire[ks348d2-1:0]  qi3b099;
wire[ks348d2-1:0]  xjc264f;
wire[ks348d2-1:0]  do993fe;
wire                    qtc9ff3;
wire                    jp4ff9d;
wire[sj2348d-1:0]  dmfe774;
wire[sj2348d-1:0]  co9dd1e;
generate         case(xj503f8)            0  :  begin                     if(wyb3750=="ADD") begin                        pmi_add #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_add"   ))                        ls83c50 (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b0       ),                           .Result     (jp6e75e          ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end else begin                        pmi_sub #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_sub"   ))                        ks92bcc (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b1       ),                           .Result     (jp6e75e          ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end                  end            1  :  begin                     if(wyb3750=="ADD") begin                        pmi_add #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_add"   ))                        ls83c50 (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b0       ),                           .Result     (pfe6b30     ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end else begin                        pmi_sub #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_sub"   ))                        ks92bcc (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b1       ),                           .Result     (pfe6b30     ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end                     lqee0f9_FFTC2048 #(.gb707ca  (1           ),                                 .mg1f2a2 (ps7340e  ))                     ir9ac93 (                           .clk  (clk     ),                           .rstn (rstn    ),                           .pfe9af9    (pfe6b30  ),                           .hdaa0f5    (jp6e75e       )                           ) ;                  end            2  :  begin                                          lqee0f9_FFTC2048 #(.gb707ca  (1              ),                                 .mg1f2a2 (sj2348d   ))                     lqd5b3a (                           .clk  (clk                         ),                           .rstn (rstn                        ),                           .pfe9af9    (ba3f16e[ps7340e-1:ks348d2]),                           .hdaa0f5    (mgacc3b                        )                           ) ;                     lqee0f9_FFTC2048 #(.gb707ca  (1              ),                                 .mg1f2a2 (sj2348d   ))                     jc52142 (                           .clk  (clk                         ),                           .rstn (rstn                        ),                           .pfe9af9    (fac5b9d[ps7340e-1:ks348d2]),                           .hdaa0f5    (ri30ec2                        )                           ) ;                     if(wyb3750=="ADD") begin                        pmi_add #( .pmi_data_width    (ks348d2  ),                                   .pmi_result_width  (ks348d2  ),                                   .pmi_sign          ("off"         ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_add"    ))                        ri867c3 (                           .DataA      (ba3f16e[ks348d2-1:0] ),                           .DataB      (fac5b9d[ks348d2-1:0] ),                           .Cin        (1'b0                ),                           .Result     (qi3b099          ),                           .Cout       (qtc9ff3            ),                           .Overflow   (                    )                        );                     end else begin                        pmi_sub #( .pmi_data_width    (ks348d2  ),                                   .pmi_result_width  (ks348d2  ),                                   .pmi_sign          ("off"         ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_sub"    ))                        wy2b883 (                           .DataA      (ba3f16e[ks348d2-1:0] ),                           .DataB      (fac5b9d[ks348d2-1:0] ),                           .Cin        (1'b1                ),                           .Result     (qi3b099          ),                           .Cout       (qtc9ff3            ),                           .Overflow   (                    )                        );                     end                     lqee0f9_FFTC2048 #(.gb707ca  (1  ),                                 .mg1f2a2 (1  ))                     rt5fa3a (                           .clk  (clk           ),                           .rstn (rstn          ),                           .pfe9af9    (qtc9ff3      ),                           .hdaa0f5    (jp4ff9d  )                           ) ;                     lqee0f9_FFTC2048 #(.gb707ca  (1              ),                                 .mg1f2a2 (ks348d2   ))                     ea5c380 (                           .clk  (clk           ),                           .rstn (rstn          ),                           .pfe9af9    (qi3b099    ),                           .hdaa0f5    (xjc264f)                           ) ;                                       lqee0f9_FFTC2048 #(.gb707ca  (1              ),                                 .mg1f2a2 (ks348d2   ))                     bl4a79a (                           .clk  (clk           ),                           .rstn (rstn          ),                           .pfe9af9    (xjc264f),                           .hdaa0f5    (do993fe )                           ) ;                     if(wyb3750=="ADD") begin                        pmi_add #( .pmi_data_width    (sj2348d ),                                   .pmi_result_width  (sj2348d ),                                   .pmi_sign          ("on"         ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_add"    ))                        nr406b0 (                           .DataA      (mgacc3b),                           .DataB      (ri30ec2),                           .Cin        (jp4ff9d                 ),                           .Result     (dmfe774                  ),                           .Cout       (                             ),                           .Overflow   (                             )                        );                     end else begin                        pmi_sub #( .pmi_data_width    (sj2348d ),
                                   .pmi_result_width  (sj2348d ),                                   .pmi_sign          ("on"         ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_sub"    ))                        uvcceb9 (                           .DataA      (mgacc3b),                           .DataB      (ri30ec2),                           .Cin        (jp4ff9d                 ),                           .Result     (dmfe774                  ),                           .Cout       (                             ),                           .Overflow   (                             )                        );                     end                     lqee0f9_FFTC2048 #(.gb707ca  (1              ),                                 .mg1f2a2 (sj2348d   ))                     mtb1c56 (                           .clk  (clk              ),                           .rstn (rstn             ),                           .pfe9af9    (dmfe774      ),                           .hdaa0f5    (co9dd1e  )                           ) ;                     assign jp6e75e = {co9dd1e,do993fe};                  end            default  :  begin                     if(wyb3750=="ADD") begin                        pmi_add #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_add"   ))                        ls83c50 (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b0       ),                           .Result     (pfe6b30     ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end else begin                        pmi_sub #( .pmi_data_width    (ps7340e  ),                                   .pmi_result_width  (ps7340e  ),                                   .pmi_sign          ("on"        ),                                   .pmi_family        (ayea07f),                                   .module_type       ("pmi_sub"   ))                        ks92bcc (                           .DataA      (ba3f16e          ),                           .DataB      (fac5b9d          ),                           .Cin        (1'b1       ),                           .Result     (pfe6b30     ),                           .Cout       (           ),                           .Overflow   (           )                        );                     end                     lqee0f9_FFTC2048 #(.gb707ca  (1           ),                                 .mg1f2a2 (ps7340e  ))                     ir9ac93 (                           .clk  (clk     ),                           .rstn (rstn    ),                           .pfe9af9    (pfe6b30  ),                           .hdaa0f5    (jp6e75e       )                           ) ;                  end         endcase      endgenerate
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module thf9cbe_FFTC2048(
               clk,            
               rstn,           
               ba3f16e,              
               fac5b9d,              
               jp6e75e,              
               pfe9af9,              
               rt6be72               
               ) ;
parameter  dzd8704 = `DATA_WIDTH+`TWID_WIDTH;
input                      clk ;
input                      rstn;
input [`DATA_WIDTH-1:0]    ba3f16e;
input [`TWID_WIDTH-1:0]    fac5b9d;
input [`DATA_WIDTH-1:0]    jp6e75e;
input [`TWID_WIDTH-1:0]    pfe9af9;
output[`DATA_WIDTH:0]    rt6be72;
wire[dzd8704:0]       alc3f66 ;
`ifdef TRUNCATE
`else
reg [`DATA_WIDTH:0]  aa1fb34;
reg                  shfd9a1;
wire ne57a3b = alc3f66[dzd8704];
`endif
`ifdef USE_MULT36
wire[dzd8704-1:0] wldcc4;
wire[dzd8704-1:0] jc7312e;
wire[dzd8704:0]   goc4b98;
wire[dzd8704:0]   ym2e60a;
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
wire[dzd8704-1:0] wldcc4;
wire[dzd8704-1:0] jc7312e;
wire[dzd8704:0]   goc4b98;
wire[dzd8704:0]   ym2e60a;
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef USE_MULT36
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef USE_MULT36
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
`endif
            
`ifdef TRUNCATE
         assign rt6be72 = {alc3f66[dzd8704],alc3f66[dzd8704-2:`TWID_WIDTH-1]};
`else
         always @(posedge clk or negedge rstn)         begin            if(!rstn) begin               aa1fb34   <= {(`DATA_WIDTH+1){1'b0}};               shfd9a1 <= 1'b0;            end else begin               aa1fb34 <= {alc3f66[dzd8704],alc3f66[dzd8704-2:`TWID_WIDTH-1]};               shfd9a1 <= ne57a3b ? (alc3f66[`TWID_WIDTH-2]&(|alc3f66[`TWID_WIDTH-3:0])) : alc3f66[`TWID_WIDTH-2];            end         end         su566ea_FFTC2048 #(.wyb3750    ("ADD"         ),                     .ps7340e (`DATA_WIDTH+1 ),                     .ayea07f (`DEVICE_FAMILY),                     .xj503f8  (1             ))         ie3e311 (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (aa1fb34   ),                  .fac5b9d       ({{`DATA_WIDTH{1'b0}},shfd9a1}),                  .jp6e75e       (rt6be72          )               );
`endif
`ifdef USE_MULT36
                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (1             ),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("DSP"         ))         hod5cd9 (                     .DataA                     (ba3f16e             ),                     .DataB                     (fac5b9d             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (wldcc4     )                  );                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (1             ),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("DSP"         ))         jcca8f5 (                     .DataA                     (jp6e75e             ),                     .DataB                     (pfe9af9             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (jc7312e     )                  );         assign goc4b98 = {wldcc4[dzd8704-1],wldcc4};         assign ym2e60a = {jc7312e[dzd8704-1],jc7312e};
                  su566ea_FFTC2048 #(.wyb3750    ("ADD"               ),                     .ps7340e (dzd8704+1        ),                     .ayea07f (`DEVICE_FAMILY),                     .xj503f8  (1+`ADDER_PIPELINE   ))         ls83c50 (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (goc4b98       ),                  .fac5b9d       (ym2e60a       ),                  .jp6e75e       (alc3f66      )               );
`endif
`ifdef HMAC_NON36
         pmi_multaddsub #( .pmi_dataa_width        (`DATA_WIDTH      ),            .pmi_datab_width        (`TWID_WIDTH      ),            .module_type            ("pmi_multaddsub" ),            .pmi_sign               ("on"             ),            .pmi_additional_pipeline(1                ),            .pmi_add_sub            ("add"            ),            .pmi_input_reg          ("on"             ),            .pmi_output_reg         ("on"             ),            .pmi_family             (`DEVICE_FAMILY   ),            .pmi_implementation     ("DSP"            ))         ls25fa2 (                           .DataA0                 (ba3f16e                ),                           .DataA1                 (jp6e75e                ),                           .DataB0                 (fac5b9d                ),                           .DataB1                 (pfe9af9                ),                           .Clock                  (clk              ),                           .ClkEn                  (1'b1             ),                           .Aclr                   (1'b0             ),                           .Result                 (alc3f66            )                        );
`endif
`ifdef DIST_MULT
                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (`MULT_PIPELINE-2),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("LUT"         ))         ie8271c (                     .DataA                     (ba3f16e             ),                     .DataB                     (fac5b9d             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (wldcc4     )                  );                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (`MULT_PIPELINE-2),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("LUT"         ))         co975fb (                     .DataA                     (jp6e75e             ),                     .DataB                     (pfe9af9             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (jc7312e     )                  );
         assign goc4b98 = {wldcc4[dzd8704-1],wldcc4};         assign ym2e60a = {jc7312e[dzd8704-1],jc7312e};
         su566ea_FFTC2048 #(.wyb3750    ("ADD"               ),                     .ps7340e (dzd8704+1        ),                     .ayea07f (`DEVICE_FAMILY),                     .xj503f8  (1+`ADDER_PIPELINE   ))         ls83c50 (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (goc4b98       ),                  .fac5b9d       (ym2e60a       ),                  .jp6e75e       (alc3f66      )               );
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module dmee6a7_FFTC2048(
               clk,            
               rstn,           
               ba3f16e,              
               fac5b9d,              
               jp6e75e,              
               pfe9af9,              
               rt6be72               
               ) ;
parameter  dzd8704 = `DATA_WIDTH+`TWID_WIDTH;
input                      clk ;
input                      rstn;
input [`DATA_WIDTH-1:0]    ba3f16e;
input [`TWID_WIDTH-1:0]    fac5b9d;
input [`DATA_WIDTH-1:0]    jp6e75e;
input [`TWID_WIDTH-1:0]    pfe9af9;
output[`DATA_WIDTH:0]    rt6be72;
wire[dzd8704:0]       alc3f66 ;
`ifdef TRUNCATE
`else
reg [`DATA_WIDTH:0]  aa1fb34;
reg                  shfd9a1;
wire ne57a3b = alc3f66[dzd8704];
`endif
`ifdef USE_MULT36
wire[dzd8704-1:0] wldcc4;
wire[dzd8704-1:0] jc7312e;
wire[dzd8704:0]   goc4b98;
wire[dzd8704:0]   ym2e60a;
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
wire[dzd8704-1:0] wldcc4;
wire[dzd8704-1:0] jc7312e;
wire[dzd8704:0]   wla4799;
wire[dzd8704:0]   tw1e66d;
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef USE_MULT36
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef USE_MULT36
`endif
`ifdef HMAC_NON36
`endif
`ifdef DIST_MULT
`endif
            
`ifdef TRUNCATE
         assign rt6be72 = {alc3f66[dzd8704],alc3f66[dzd8704-2:`TWID_WIDTH-1]};
`else
         always @(posedge clk or negedge rstn)         begin            if(!rstn) begin               aa1fb34   <= {(`DATA_WIDTH+1){1'b0}};               shfd9a1 <= 1'b0;            end else begin               aa1fb34 <= {alc3f66[dzd8704],alc3f66[dzd8704-2:`TWID_WIDTH-1]};               shfd9a1 <= ne57a3b ? (alc3f66[`TWID_WIDTH-2]&(|alc3f66[`TWID_WIDTH-3:0])) : alc3f66[`TWID_WIDTH-2];            end         end         su566ea_FFTC2048 #(.wyb3750    ("ADD"         ),                     .ps7340e (`DATA_WIDTH+1 ),                     .xj503f8  (1             ))         ie3e311 (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (aa1fb34   ),                  .fac5b9d       ({{`DATA_WIDTH{1'b0}},shfd9a1} ),                  .jp6e75e       (rt6be72          )               );
`endif
`ifdef USE_MULT36
                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (1             ),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("DSP"         ))         hod5cd9 (                     .DataA                     (ba3f16e             ),                     .DataB                     (fac5b9d             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (wldcc4     )                  );                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (1             ),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("DSP"         ))         jcca8f5 (                     .DataA                     (jp6e75e             ),                     .DataB                     (pfe9af9             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (jc7312e     )                  );         assign goc4b98 = {wldcc4[dzd8704-1],wldcc4};         assign ym2e60a = {jc7312e[dzd8704-1],jc7312e};
                  su566ea_FFTC2048 #(.wyb3750    ("SUB"               ),                     .ps7340e (dzd8704+1        ),                     .ayea07f (`DEVICE_FAMILY),                     .xj503f8  (1+`ADDER_PIPELINE   ))         ls83c50 (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (goc4b98       ),                  .fac5b9d       (ym2e60a       ),                  .jp6e75e       (alc3f66      )               );
`endif
`ifdef HMAC_NON36
         pmi_multaddsub #( .pmi_dataa_width        (`DATA_WIDTH      ),            .pmi_datab_width        (`TWID_WIDTH      ),            .module_type            ("pmi_multaddsub" ),            .pmi_sign               ("on"             ),            .pmi_additional_pipeline(1                ),            .pmi_add_sub            ("sub"            ),            .pmi_input_reg          ("on"             ),            .pmi_output_reg         ("on"             ),            .pmi_family             (`DEVICE_FAMILY   ),            .pmi_implementation     ("DSP"            ))         ls25fa2 (                           .DataA0                 (ba3f16e                ),                           .DataA1                 (jp6e75e                ),                           .DataB0                 (fac5b9d                ),                           .DataB1                 (pfe9af9                ),                           .Clock                  (clk              ),                           .ClkEn                  (1'b1             ),                           .Aclr                   (1'b0             ),                           .Result                 (alc3f66            )                        );
`endif
`ifdef DIST_MULT
                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (`MULT_PIPELINE-2),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("LUT"         ))         ie8271c (                     .DataA                     (ba3f16e             ),                     .DataB                     (fac5b9d             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (wldcc4     )                  );                  pmi_mult #( .pmi_dataa_width           (`DATA_WIDTH   ),      .pmi_datab_width           (`TWID_WIDTH   ),      .module_type               ("pmi_mult"    ),      .pmi_sign                  ("on"          ),      .pmi_additional_pipeline   (`MULT_PIPELINE-2),      .pmi_input_reg             ("on"          ),      .pmi_output_reg            ("on"          ),      .pmi_family                (`DEVICE_FAMILY),      .pmi_implementation        ("LUT"         ))         co975fb (                     .DataA                     (jp6e75e             ),                     .DataB                     (pfe9af9             ),                     .Clock                     (clk           ),                     .ClkEn                     (1'b1          ),                     .Aclr                      (1'b0          ),                     .Result                    (jc7312e     )                  );
         assign wla4799 = {wldcc4[dzd8704-1],wldcc4};         assign tw1e66d = {jc7312e[dzd8704-1],jc7312e};         su566ea_FFTC2048 #(.wyb3750    ("SUB"               ),                     .ps7340e (dzd8704+1        ),                     .ayea07f (`DEVICE_FAMILY),                     .xj503f8  (1+`ADDER_PIPELINE   ))         ks92bcc (                  .rstn    (rstn       ),                  .clk     (clk        ),                  .ba3f16e       (wla4799       ),                  .fac5b9d       (tw1e66d       ),                  .jp6e75e       (alc3f66      )               );
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module lqee0f9_FFTC2048(
             rstn,                  
             clk,                   
             pfe9af9,                     
             hdaa0f5                      
             ) ;
parameter      gb707ca  = 3;
parameter      mg1f2a2 = 16;
input                   rstn;
input                   clk;
input [mg1f2a2-1:0]   pfe9af9;
output[mg1f2a2-1:0]   hdaa0f5;
reg [mg1f2a2-1:0]     yz95d45[0:gb707ca-1];
integer                 en75165;
always @(posedge clk or negedge rstn)      begin         if(!rstn)            for(en75165=0;en75165<gb707ca;en75165=en75165+1) yz95d45[en75165] <= {mg1f2a2{1'b0}};         else begin            yz95d45[0] <= pfe9af9;            for(en75165=1;en75165<gb707ca;en75165=en75165+1) yz95d45[en75165] <= yz95d45[en75165-1];         end      end
      assign hdaa0f5 = yz95d45[gb707ca-1];
   endmodule                                                                                       
`ifdef BFPU_PRESENT
`timescale 1 ns / 100 ps
module tw3016e_FFTC2048 (
                  rstn,                
                  clk,                 
                  rv2dca9,               
                  dz6e54e,               
                  su72a76,               
                  oh953b0,               
               `ifdef BFPU_PRESENT
                  uka9d85,
                  al4ec28,              
                  fa76144,
                  tjb0a23,                
               `ifdef BIT_REVERSE
                  an8511f,
               `endif
                  db288fc,              
                  uv447e6,              
                  exponent,            
                  qi1f9a5,
                  cz709f8,
                  ibend,
               `endif
                  ks34a7f,               
                  hda53f9,               
                  an29fcf,               
                  xj4fe7c                
               ) ;
parameter   ip7f3e6 = `WR_LATENCY+2;
input                   rstn;
input                   clk;
input [`DATA_WIDTH+1:0] rv2dca9;
input [`DATA_WIDTH+1:0] dz6e54e;
input [`DATA_WIDTH+1:0] su72a76;
input [`DATA_WIDTH+1:0] oh953b0;
`ifdef BFPU_PRESENT
input                   uka9d85;
input                   fa76144;
input                   al4ec28;
input [`LOG2_NBY2-1:0]  tjb0a23;
`ifdef BIT_REVERSE
input [`LOG2_NBY2-1:0]  an8511f;
`endif
input [`LOG2_NBY2-1:0]  db288fc;
input                   qi1f9a5;
input                   ibend;
input                   uv447e6;
output[1:0]             cz709f8;
output[`STAGE_WIDTH:0]  exponent;
`endif
output[`DATA_WIDTH+1:0] ks34a7f;
output[`DATA_WIDTH+1:0] hda53f9;
output[`DATA_WIDTH+1:0] an29fcf;
output[`DATA_WIDTH+1:0] xj4fe7c;
reg [`DATA_WIDTH+1:0]   ks34a7f;
reg [`DATA_WIDTH+1:0]   hda53f9;
reg [`DATA_WIDTH+1:0]   an29fcf;
reg [`DATA_WIDTH+1:0]   xj4fe7c;
reg [`DATA_WIDTH+1:0]   ohd391;
reg [`DATA_WIDTH+1:0]   ne69c8c;
reg [`DATA_WIDTH+1:0]   wj4e462;
reg [`DATA_WIDTH+1:0]   cm72315;
reg [`DATA_WIDTH+1:0]   vx918a9;
reg [`DATA_WIDTH+1:0]   vk8c54e;
reg [`DATA_WIDTH+1:0]   qg62a72;
reg [`DATA_WIDTH+1:0]   sw15391;
`ifdef BFPU_PRESENT
reg [1:0]               cz709f8;
reg [`STAGE_WIDTH:0]    wj4e448;
reg [`STAGE_WIDTH:0]    exponent;
reg [ip7f3e6-1:0]    zm8914f;
`endif
wire                    xw48a7a;
wire                    nr453d3;
reg [1:0]               cb29e9e;
reg [`LOG2_NBY2-1:0]    nr4f4f4;
reg [`LOG2_NBY2-1:0]    kd7a7a7;
reg [1:0]               kdd3d3d;
wire[`LOG2_NBY2-1:0]    rv9e9ed;
reg [1:0]               xwf4f6f;
reg [`LOG2_NBY2-1:0]    fca7b7b;
reg [`LOG2_NBY2-1:0]    lf3dbdb;
wire[1:0]               shededf;
reg [`LOG2_NBY2-1:0]    kd6f6fc;
wire                    zx7b7e4;
wire                    ykdbf27;
integer                 en75165;
`ifdef BFPU_PRESENT
wire                 blfc9cb;
wire[`LOG2_NBY2-1:0] pse4e5f;
reg [`LOG2_NBY2-1:0] jr272fa[ip7f3e6-1:0];
`ifdef TRUNCATE
wire[`LOG2_NBY2-1:0] uicbeb4 = jr272fa[ip7f3e6-3];
`else
wire[`LOG2_NBY2-1:0] uicbeb4 = jr272fa[ip7f3e6-4];
`endif
reg                  db6166;
reg                  do30b37;
reg [1:0]            cb859bb;
reg [1:0]            wl2cddd;
reg [1:0]            ps66eec;
reg [1:0]            nt37763;
reg [`LOG2_NBY2-1:0] epbbb1f;
reg [`LOG2_NBY2-1:0] lddd8fc[0:ip7f3e6];
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BIT_REVERSE
reg [`LOG2_NBY2-1:0] rg63f37;
`endif
`ifdef TRUNCATE
`ifdef BIT_REVERSE
`else
`endif
`else
`ifdef BIT_REVERSE
`else
`endif
`endif
`endif
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BIT_REVERSE
`endif
`ifdef TRUNCATE
`ifdef BIT_REVERSE
`else
`endif
`else
`ifdef BIT_REVERSE
`else
`endif
`endif
`endif
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BIT_REVERSE
`endif
`ifdef TRUNCATE
`ifdef BIT_REVERSE
`else
`endif
`else
`ifdef BIT_REVERSE
`else
`endif
`endif
`endif
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`ifdef BFPU_PRESENT
`endif
      
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ohd391  <= {(`DATA_WIDTH+2){1'b0}};            ne69c8c  <= {(`DATA_WIDTH+2){1'b0}};            wj4e462  <= {(`DATA_WIDTH+2){1'b0}};            cm72315  <= {(`DATA_WIDTH+2){1'b0}};            vx918a9 <= {(`DATA_WIDTH+2){1'b0}};            vk8c54e <= {(`DATA_WIDTH+2){1'b0}};            qg62a72 <= {(`DATA_WIDTH+2){1'b0}};            sw15391 <= {(`DATA_WIDTH+2){1'b0}};            ks34a7f    <= {(`DATA_WIDTH+2){1'b0}};            hda53f9    <= {(`DATA_WIDTH+2){1'b0}};            an29fcf    <= {(`DATA_WIDTH+2){1'b0}};            xj4fe7c    <= {(`DATA_WIDTH+2){1'b0}};         end else begin            ohd391  <= rv2dca9;            ne69c8c  <= dz6e54e;            wj4e462  <= su72a76;            cm72315  <= oh953b0;            vx918a9 <= ohd391;            vk8c54e <= ne69c8c;            qg62a72 <= wj4e462;            sw15391 <= cm72315;            ks34a7f    <= vx918a9;            hda53f9    <= vk8c54e;            an29fcf    <= qg62a72;            xj4fe7c    <= sw15391;         end      end
`ifdef BFPU_PRESENT
`ifdef TRUNCATE
`else
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            for(en75165=0;en75165<ip7f3e6;en75165=en75165+1) lddd8fc[en75165] <= {`LOG2_NBY2{1'b0}};         else begin            lddd8fc[0] <= db288fc;            for(en75165=1;en75165<ip7f3e6;en75165=en75165+1) lddd8fc[en75165] <= lddd8fc[en75165-1];         end      end
`ifdef TRUNCATE
      assign blfc9cb = zm8914f[ip7f3e6-5];      assign zx7b7e4   = zm8914f[ip7f3e6-6];      assign ykdbf27     = rv9e9ed==lddd8fc[ip7f3e6-8];
`else
      assign blfc9cb = zm8914f[ip7f3e6-6];      assign zx7b7e4   = zm8914f[ip7f3e6-7];      assign ykdbf27     = rv9e9ed==lddd8fc[ip7f3e6-9];
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) zm8914f <= {ip7f3e6{1'b0}};         else      zm8914f <= {zm8914f[ip7f3e6-2:0],al4ec28};      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn)            for(en75165=0;en75165<ip7f3e6;en75165=en75165+1) jr272fa[en75165] <= {`LOG2_NBY2{1'b0}};         else begin            jr272fa[0] <= tjb0a23;            for(en75165=1;en75165<ip7f3e6;en75165=en75165+1) jr272fa[en75165] <= jr272fa[en75165-1];         end      end
      
`ifdef TRUNCATE
      assign rv9e9ed     = jr272fa[ip7f3e6-6];      assign pse4e5f = jr272fa[ip7f3e6-5];
`else
      assign rv9e9ed     = jr272fa[ip7f3e6-7];      assign pse4e5f = jr272fa[ip7f3e6-6];
`endif
`ifdef BIT_REVERSE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            rg63f37 <= {`LOG2_NBY2{1'b0}};         else for(en75165=0;en75165<`LOG2_NBY2;en75165=en75165+1)            rg63f37[en75165] <= an8511f[`LOG2_NBY2-1-en75165];      end
`endif
   
`ifdef TRUNCATE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            kd6f6fc <= 0;         else
`ifdef BIT_REVERSE
            kd6f6fc <= fa76144 ? rg63f37 :                        {jr272fa[ip7f3e6-8][`LOG2_NBY2-2:0],jr272fa[ip7f3e6-8][`LOG2_NBY2-1]};
`else
            kd6f6fc <= fa76144 ? jr272fa[1] :                        {jr272fa[ip7f3e6-8][`LOG2_NBY2-2:0],jr272fa[ip7f3e6-8][`LOG2_NBY2-1]};
`endif
      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            kd6f6fc <= 0;         else
`ifdef BIT_REVERSE
            kd6f6fc <= fa76144 ? rg63f37 :                        {jr272fa[ip7f3e6-9][`LOG2_NBY2-2:0],jr272fa[ip7f3e6-9][`LOG2_NBY2-1]};
`else
            kd6f6fc <= fa76144 ? jr272fa[1] :                        {jr272fa[ip7f3e6-9][`LOG2_NBY2-2:0],jr272fa[ip7f3e6-9][`LOG2_NBY2-1]};
`endif
      end
`endif
            assign xw48a7a = ((|rv2dca9[`DATA_WIDTH+1:`DATA_WIDTH])&(!(&rv2dca9[`DATA_WIDTH+1:`DATA_WIDTH]))) ||                      ((|dz6e54e[`DATA_WIDTH+1:`DATA_WIDTH])&(!(&dz6e54e[`DATA_WIDTH+1:`DATA_WIDTH]))) ||                      ((|su72a76[`DATA_WIDTH+1:`DATA_WIDTH])&(!(&su72a76[`DATA_WIDTH+1:`DATA_WIDTH]))) ||                      ((|oh953b0[`DATA_WIDTH+1:`DATA_WIDTH])&(!(&oh953b0[`DATA_WIDTH+1:`DATA_WIDTH])));      assign nr453d3 = ((|rv2dca9[`DATA_WIDTH+1:`DATA_WIDTH-1])&(!(&rv2dca9[`DATA_WIDTH+1:`DATA_WIDTH-1]))) ||                      ((|dz6e54e[`DATA_WIDTH+1:`DATA_WIDTH-1])&(!(&dz6e54e[`DATA_WIDTH+1:`DATA_WIDTH-1]))) ||                      ((|su72a76[`DATA_WIDTH+1:`DATA_WIDTH-1])&(!(&su72a76[`DATA_WIDTH+1:`DATA_WIDTH-1]))) ||                      ((|oh953b0[`DATA_WIDTH+1:`DATA_WIDTH-1])&(!(&oh953b0[`DATA_WIDTH+1:`DATA_WIDTH-1])));
      always @(posedge clk or negedge rstn)      begin         if(!rstn)               db6166 <= 1'b0;         else if(ykdbf27 && fa76144) db6166 <= 1'b1;         else if(db6166 && ykdbf27)    db6166 <= 1'b0;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            do30b37 <= 1'b0;         else if(db6166 && ykdbf27) do30b37 <= 1'b1;         else                 do30b37 <= 1'b0;      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            xwf4f6f   <= 2'b00;            fca7b7b <= {`LOG2_NBY2{1'b0}};            lf3dbdb <= {`LOG2_NBY2{1'b0}};         end else if(do30b37 || ibend) begin            xwf4f6f   <= 2'b00;            fca7b7b <= {`LOG2_NBY2{1'b0}};            lf3dbdb <= {`LOG2_NBY2{1'b0}};         end else if(ykdbf27 && zx7b7e4) begin            case({xw48a7a,nr453d3})               2'b01 :  begin                           lf3dbdb <= kd7a7a7;                           if(cb29e9e==2'b00) begin                              xwf4f6f <= 2'b01;                              if(uka9d85) fca7b7b <= pse4e5f;                              else             fca7b7b <= rv9e9ed;                           end else begin                              xwf4f6f   <= cb29e9e;                              fca7b7b <= nr4f4f4;                           end                        end               2'b11 :  begin                           fca7b7b <= nr4f4f4;                           xwf4f6f <= 2'b11;                           if(cb29e9e!=2'b11) begin                              if(uka9d85) lf3dbdb <= pse4e5f;                              else             lf3dbdb <= rv9e9ed;                           end else begin                              lf3dbdb <= kd7a7a7;                           end                        end               default: begin                           xwf4f6f   <= cb29e9e;                           fca7b7b <= nr4f4f4;                           lf3dbdb <= kd7a7a7;                        end            endcase         end      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn)            cb859bb <= 2'b00;         else if(do30b37 || ibend)            cb859bb <= 2'b00;         else if(ykdbf27 && zx7b7e4)            case({xw48a7a,nr453d3})               2'b00 :  if(!(kd7a7a7==0))      cb859bb <= 2'b10;                        else if(!(nr4f4f4==0)) cb859bb <= 2'b01;                        else                  cb859bb <= 2'b00;               2'b01 :  if(!(kd7a7a7==0))      cb859bb <= 2'b10;                        else if(!(nr4f4f4==0)) cb859bb <= 2'b01;                        else if(cz709f8==0)     cb859bb <= 2'b01;                        else                  cb859bb <= 2'b00;               2'b10,               2'b11 :  if(!(kd7a7a7==0))      cb859bb <= 2'b10;                        else if(cz709f8==2'b00) cb859bb <= 2'b10;                        else if(cz709f8==2'b01) cb859bb <= 2'b01;                        else if(!(nr4f4f4==0)) cb859bb <= 2'b01;                        else                  cb859bb <= 2'b00;            endcase      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn)            wl2cddd <= 2'b00;         else casex(xwf4f6f)            2'b00 :  wl2cddd <= 2'b00;            2'b01 :  if(kd6f6fc < fca7b7b)      wl2cddd <= 2'b01;                     else                      wl2cddd <= 2'b00;            2'b1x :  if(kd6f6fc < fca7b7b)      wl2cddd <= 2'b10;                     else if(kd6f6fc < lf3dbdb) wl2cddd <= 2'b01;                     else                      wl2cddd <= 2'b00;         endcase      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            epbbb1f <= 0;         else            epbbb1f <= kd6f6fc;      end
                assign shededf = qi1f9a5==1 ? wl2cddd : epbbb1f==0 ? cb859bb : wl2cddd;   
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            cb29e9e      <= 2'b00;            nr4f4f4    <= {`LOG2_NBY2{1'b0}};            kd7a7a7    <= {`LOG2_NBY2{1'b0}};            ps66eec <= 2'b00;         end else if(do30b37 || ibend) begin            cb29e9e      <= 2'b00;            nr4f4f4    <= {`LOG2_NBY2{1'b0}};            kd7a7a7    <= {`LOG2_NBY2{1'b0}};            ps66eec <= 2'b00;         end else case({xw48a7a,nr453d3,shededf})               4'b0100,               4'b1101  :  if(cb29e9e==2'b00) begin                              cb29e9e   <= 2'b01;                              if(uka9d85) begin                                 nr4f4f4 <= pse4e5f;                                 ps66eec <= 2'b01;                              end else begin                                 nr4f4f4 <= rv9e9ed;                                 ps66eec <= 2'b00;                              end                           end else ps66eec <= 2'b00;               4'b1100  :  begin                              cb29e9e   <= 2'b11;                              if(cb29e9e!=2'b11) begin                                 if(uka9d85) begin                                    kd7a7a7 <= pse4e5f;                                    ps66eec <= 2'b10;                                 end else begin                                    kd7a7a7 <= rv9e9ed;                                    ps66eec <= 2'b00;                                 end                              end else ps66eec <= 2'b00;                           end               default  :  begin                              if(rv9e9ed==0) begin                                 cb29e9e   <= 2'b00;                                 nr4f4f4 <= {`LOG2_NBY2{1'b0}};                                 kd7a7a7 <= {`LOG2_NBY2{1'b0}};                              end                              ps66eec <= 2'b00;                           end            endcase      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) nt37763 <= 2'b00;         else      nt37763 <= shededf;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) kdd3d3d <= 2'b00;         else casex({cb29e9e,nt37763})            4'b0101,            4'bxx10,            4'b11xx  :  kdd3d3d <= 2'b10;            4'b0001,            4'b0100  :  kdd3d3d <= 2'b01;            default  :  kdd3d3d <= 2'b00;         endcase      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)          cz709f8 <= 2'b00;         else if(qi1f9a5) cz709f8 <= shededf;         else               cz709f8 <= kdd3d3d + ps66eec;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            wj4e448 <= 0;         else if(do30b37 || ibend)            wj4e448 <= 0;         else if(uicbeb4==db288fc && zm8914f[ip7f3e6-2])            wj4e448 <= wj4e448 + cz709f8;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            exponent <= 0;         else if(uv447e6)            exponent <= wj4e448;         else            exponent <= 0;      end
`endif
   endmodule
`endif
                                                                                          
`timescale 1 ns / 100 ps
module sj12f6f_FFTC2048 (
              clk,               
              rstn,              
              fft_mode,          
              dire,              
              diim,              
              dore,              
              doim               
              ) ;
input                      clk;
input                      rstn;
input                      fft_mode ;
input [`DATA_WIDTH-1:0]    dire;
input [`DATA_WIDTH-1:0]    diim;
output [`DATA_WIDTH-1:0]    dore;
output [`DATA_WIDTH-1:0]    doim;
reg [`DATA_WIDTH-1:0]      dore;
reg [`DATA_WIDTH-1:0]      doim;
                        always @(posedge clk or negedge rstn)      begin         if(!rstn)            doim <= {`DATA_WIDTH{1'b0}};         else            doim <= fft_mode ? (1'b1 + (~diim)) : diim;      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) dore <= {`DATA_WIDTH{1'b0}};         else      dore <= dire;      end
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module jpc7848_FFTC2048 (
               clk,                 
               rstn,                
            `ifdef DYNAMIC_POINTS
               points,              
               xw48d1e,          
            `endif
            `ifdef MODE_PORT_READ
               mode,                
               co34798,            
            `endif
            `ifdef SFACT_PORT_READ
               sfact,               
               do1e601,           
            `endif
               nrf300a,            
               co98057,               
               hoc02b9,               
            `ifdef DYNAMIC_POINTS
               fc15ca,            
               ouae52,        
            `endif
            `ifdef MODE_PORT_READ
               ne57290,              
               ieb9482,          
            `endif
            `ifdef SFACT_PORT_READ
               psca410,             
               zk52083,         
            `endif
               cb9041a,          
               co820d5,             
               uk106a9              
               );
input                       clk;
input                       rstn;
`ifdef DYNAMIC_POINTS
input [`NFFT_WIDTH-1:0]     points;
input                       xw48d1e;
`endif
`ifdef MODE_PORT_READ
input                       mode;
input                       co34798;
`endif
`ifdef SFACT_PORT_READ
input [`SFACT_WIDTH-1:0]    sfact;
input                       do1e601;
`endif
input                       nrf300a;
input [`DIN_WIDTH-1:0]     co98057;
input [`DIN_WIDTH-1:0]     hoc02b9;
`ifdef DYNAMIC_POINTS
output[`NFFT_WIDTH-1:0]     fc15ca;
output                      ouae52;
`endif
`ifdef MODE_PORT_READ
output                      ne57290;
output                      ieb9482;
`endif
`ifdef SFACT_PORT_READ
output[`SFACT_WIDTH-1:0]    psca410;
output                      zk52083;
`endif
output                      cb9041a;
output[`DIN_WIDTH-1:0]     co820d5;
output[`DIN_WIDTH-1:0]     uk106a9;
`ifdef DYNAMIC_POINTS
reg [`NFFT_WIDTH-1:0]       fc15ca;
reg                         ouae52;
`endif
`ifdef MODE_PORT_READ
reg                         ne57290;
reg                         ieb9482;
`endif
`ifdef SFACT_PORT_READ
reg [`SFACT_WIDTH-1:0]      psca410;
reg                         zk52083;
`endif
reg                         cb9041a;
reg [`DIN_WIDTH-1:0]       co820d5;
reg [`DIN_WIDTH-1:0]       uk106a9;
reg [`DIN_WIDTH-1:0]       twa83a5;
reg [`DIN_WIDTH-1:0]       wj41d2b;
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
      
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
      
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
      
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin
`ifdef DYNAMIC_POINTS
            fc15ca   <= {`NFFT_WIDTH{1'b1}};            ouae52 <= 1'b0;
`endif
`ifdef MODE_PORT_READ
            ne57290     <= 1'b0;            ieb9482 <= 1'b0;
`endif
`ifdef SFACT_PORT_READ
            psca410     <= {`SFACT_WIDTH{1'b0}};            zk52083 <= 1'b0;
`endif
            cb9041a <= 1'b0;            co820d5    <= {`DIN_WIDTH{1'b0}};            uk106a9    <= {`DIN_WIDTH{1'b0}};            twa83a5     <= {`DIN_WIDTH{1'b0}};            wj41d2b     <= {`DIN_WIDTH{1'b0}};         end else begin
`ifdef DYNAMIC_POINTS
            fc15ca     <= points;            ouae52 <= xw48d1e;
`endif
`ifdef MODE_PORT_READ
            ne57290     <= mode;            ieb9482 <= co34798;
`endif
`ifdef SFACT_PORT_READ
            psca410     <= sfact;            zk52083 <= do1e601;
`endif
            cb9041a <= nrf300a;            co820d5    <= twa83a5;            uk106a9    <= wj41d2b;            twa83a5     <= co98057;            wj41d2b     <= hoc02b9;         end      end
   endmodule                                                                                                   
`timescale 1 ns / 100 ps
module ymb9ff3_FFTC2048 (
                  rstn,                
                  clk,                 
                  vife654,         
               `ifdef DYNAMIC_POINTS
                  points,              
                  pu9951f,           
               `endif
               `ifdef MODE_PORT_READ
                  mode,                
                  modeset,             
               `endif
               `ifdef SFACT_PORT_READ
                  sfact,               
                  sfactset,            
               `endif
               `ifdef BFPU_PRESENT
               `else
               `ifdef SFACT_UNSCALE
               `else
                  dmfb548,             
               `endif
               `endif
                  jc52b77,           
                  ir95bbb,           
               `ifdef BFPU_PRESENT
               `else
                  aaacedc,              
               `endif
   
               `ifdef BFPU_PRESENT
                  uka9d85,
                  al4ec28,
                  fa76144,
                  qi1f9a5,
                  uvd9450,
               `endif
                  vica285,            
                  wj5142b,             
                  ir8a15d,             
                  xj50aed,           
                  mt8576e,             
                  sw2bb74,
                  ne5dba1,
                  db288fc,
                  fn6e854,
   
                  pf742a7,               
                  qva153e,               
                  tjb0a23,                
                  uv54fa8,              
                  nga7d44,              
                  uk3ea23,                
                  gof5118,                
                  vka88c0,            
                  ip44602,            
                  oh23014,           
   
                  rfib,                
                  ibend,               
               `ifdef BFPU_PRESENT
               `else
               `ifdef SFACT_UNSCALE
               `else
                  except,              
               `endif
               `endif
   
   
               `ifdef OUTVALID_SEL
                  ng14954,              
                                       
               `endif
   
                  obstart,             
                  outvalid             
               );
parameter   ri2a8a3 = `WR_LATENCY>8 ? `WR_LATENCY : 9;
`ifdef BIT_REVERSE
parameter   gb5451b     = 5'h01;
parameter   jea28dd    = 5'h02;
parameter   pu146eb    = 5'h04;
parameter   coa375b     = 5'h08;
parameter   hq1bad8     = 5'h10;
`else
parameter   gb5451b     = 7'h01;
parameter   jea28dd    = 7'h02;
parameter   pu146eb    = 7'h04;
parameter   coa375b     = 7'h08;
parameter   hq1bad8     = 7'h10;
parameter   ym1f53c  = 7'h20;
parameter   wwfa9e0  = 7'h40;
`endif
input                      rstn;
input                      clk;
input                      vife654;
`ifdef DYNAMIC_POINTS
input [`NFFT_WIDTH-1:0]    points;
input                      pu9951f;
`endif
`ifdef MODE_PORT_READ
input                      mode;
input                      modeset;
`endif
`ifdef SFACT_PORT_READ
input [`SFACT_WIDTH-1:0]   sfact;
input                      sfactset;
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
input                      dmfb548;
`endif
`endif
output                     jc52b77;
output                     ir95bbb;
`ifdef BFPU_PRESENT
`else
output[1:0]                aaacedc;
`endif
`ifdef BFPU_PRESENT
output                     al4ec28;
output                     fa76144;
output                     uka9d85;
output                     qi1f9a5;
output                     uvd9450;
`endif
output                     vica285;
output                     wj5142b;
output                     ir8a15d;
output                     xj50aed;
output                     mt8576e;
output[`LOG2_N-6:0]        sw2bb74;
output[`STAGE_WIDTH-1:0]   ne5dba1;
output[`LOG2_NBY2-1:0]     db288fc;
output[3:0]                fn6e854;
output                     pf742a7;
output                     qva153e;
output[`LOG2_NBY2-1:0]     tjb0a23;
output[`STAGE_WIDTH-1:0]   uv54fa8;
output[`STAGE_WIDTH-1:0]   nga7d44;
output                     uk3ea23;
output                     gof5118;
output                     vka88c0;
output                     ip44602;
output                     oh23014;
output                     rfib;
output                     ibend;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
output                     except;
`endif
`endif
`ifdef OUTVALID_SEL
output                     ng14954;
`endif
output                     obstart;
output                     outvalid;
reg                        uka9d85;
reg [`LOG2_NBY2-1:0]       tjb0a23;
reg [`LOG2_NBY2-1:0]       kq5394e;
reg [`STAGE_WIDTH-1:0]     uv54fa8;
reg [`STAGE_WIDTH-1:0]     nga7d44;
wire                       xj50aed;
integer                    en75165;
wire                       ibstart;
reg                        rfib;
reg [ri2a8a3-1:0]         uv447e6;
reg [`WR_LATENCY-1:0]      al65d63;
wire                       qi2eb1c;
wire                       yx758e1;
wire                       mgac70d;
reg                        rg63869;
reg                        db1c34b;
reg                        vka88c0,ip44602;
reg                        rg697d4,gb4bea3;
reg                        dz5f51c;
reg [`WR_LATENCY:0]        kqfa8e6;
reg                        pf742a7;
reg [`WR_LATENCY+1:0]      swa3981;
reg                        uk3ea23;
reg                        obstart;
reg [7:0]                  je30276;
`ifdef BIT_REVERSE
reg [4:0]                  vx813b2,ph9d96;
`else
reg [6:0]                  vx813b2,ph9d96;
`endif
`ifdef DYNAMIC_POINTS
reg [`LOG2_N-6:0]       sw2bb74;
reg [`LOG2_NBY2-1:0]    db288fc;
reg [`STAGE_WIDTH-1:0]  ne5dba1;
reg [3:0]               fn6e854;
reg [`NFFT_WIDTH-1:0]   ne73079;
reg [`NFFT_WIDTH-1:0]   ym1a686;
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`else
wire[`LOG2_N-6:0]       sw2bb74;
wire[3:0]               fn6e854;
wire[`LOG2_NBY2-1:0]    db288fc;
wire[`STAGE_WIDTH-1:0]  ne5dba1;
`endif
`ifdef MODE_PORT_READ
reg                           tu7c95b;
reg                           rv8489b;
reg                           ir95bbb;
reg                           jc52b77;
`else
`ifdef MODE_FORWARD
`else
`endif
`endif
`ifdef SFACT_PORT_READ
reg [`SFACT_WIDTH-1:0]     lf137ce;
reg [`SFACT_WIDTH-1:0]     ri9c793;
`else
wire[`SFACT_WIDTH-1:0]  lf137ce = {`SFACT_WIDTH{1'b0}};
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
reg   nrf9dba;
`else
`endif
`ifdef BIT_REVERSE
`ifdef DYNAMIC_POINTS
`else
`endif
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef OUTVALID_SEL
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
reg   ibend;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
reg         by76eb8;
reg         except;
`ifdef SFACT_PORT_READ
reg [1:0]   aaacedc;
reg [1:0]   cz709f8;
reg [1:0]   bab84f6[0:`WR_LATENCY-1];
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef SFACT_UNSCALE
wire[1:0]   aaacedc = 2'b00;
`endif
`ifdef SFACT_RS111
reg[1:0]    aaacedc;
`endif
`ifdef SFACT_RS211
reg [1:0]   aaacedc;
reg [`WR_LATENCY-1:0]   pff65ff;
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef DYNAMIC_POINTS
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`else
`endif
`ifdef MODE_PORT_READ
`else
`ifdef MODE_FORWARD
`else
`endif
`endif
`ifdef SFACT_PORT_READ
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`ifdef DYNAMIC_POINTS
`else
`endif
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef OUTVALID_SEL
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`ifdef SFACT_PORT_READ
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef SFACT_UNSCALE
`endif
`ifdef SFACT_RS111
`endif
`ifdef SFACT_RS211
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef DYNAMIC_POINTS
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`else
`endif
`ifdef MODE_PORT_READ
`else
`ifdef MODE_FORWARD
`else
`endif
`endif
`ifdef SFACT_PORT_READ
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef BIT_REVERSE
`ifdef DYNAMIC_POINTS
`else
`endif
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef OUTVALID_SEL
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`ifdef SFACT_PORT_READ
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef SFACT_UNSCALE
`endif
`ifdef SFACT_RS111
`endif
`ifdef SFACT_RS211
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`endif
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
      
`ifdef OUTVALID_SEL
`endif
   
`ifdef BIT_REVERSE
`else
`endif
      assign ibstart = vife654 && rfib;
      
`ifdef DYNAMIC_POINTS
`ifdef BIT_REVERSE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ne73079 <= `LOG2_N;         else if(pu9951f && !outvalid) begin            if(points < 6)       ne73079 <= 6;            else if(points > 14) ne73079 <= 14;            else                 ne73079 <= points;         end      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ne73079 <= `LOG2_N;         else if(pu9951f) begin            if(points < 6)       ne73079 <= 6;            else if(points > 14) ne73079 <= 14;            else                 ne73079 <= points;         end      end
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ym1a686 <= {`NFFT_WIDTH{1'b0}};         else      ym1a686 <= ne73079 - 1;      end
`ifdef BIT_REVERSE
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            sw2bb74   <= 1'b1;            fn6e854   <= 4'h0;            ne5dba1 <= `NUM_STAGES-1;         end else if(ibstart) begin            if(pu9951f && !outvalid) begin               sw2bb74   <= 1 << (`NUM_STAGES-points);               fn6e854   <= (`NUM_STAGES-points);               ne5dba1 <= points - 1'b1;            end else begin               sw2bb74   <= 1 << (`NUM_STAGES-ne73079);               fn6e854   <= (`NUM_STAGES-ne73079);               ne5dba1 <= ne73079 - 1'b1;            end         end      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            sw2bb74   <= 1'b1;            fn6e854   <= 4'h0;            ne5dba1 <= `NUM_STAGES-1;         end else if(ibstart) begin            if(pu9951f) begin               sw2bb74   <= 1 << (`NUM_STAGES-points);               fn6e854   <= (`NUM_STAGES-points);               ne5dba1 <= points - 1'b1;            end else begin               sw2bb74   <= 1 << (`NUM_STAGES-ne73079);               fn6e854   <= (`NUM_STAGES-ne73079);               ne5dba1 <= ne73079 - 1'b1;            end         end      end
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) db288fc <= {`LOG2_N{1'b1}};         else      db288fc <= `NUM_POINTS/2 - sw2bb74;      end
`else
      assign sw2bb74   = 1'b1;      assign fn6e854   = 4'h0;      assign db288fc   = `NUM_POINTS/2 - 1'b1;      assign ne5dba1 = `NUM_STAGES - 1'b1;
`endif
      
`ifdef MODE_PORT_READ
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            tu7c95b <= 1'b0;            rv8489b <= 1'b0;         end else begin            if(modeset)  tu7c95b <= mode;            if(ibstart) begin               if(modeset) rv8489b <= mode;               else        rv8489b <= tu7c95b;            end         end      end            always @(posedge clk or negedge rstn)      begin         if(!rstn)                 ir95bbb <= 1'b0;         else if(uv54fa8>=ne5dba1) ir95bbb <= rv8489b;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) jc52b77 <= 1'b0;         else      jc52b77 <= ibstart ? (modeset ? mode : tu7c95b) : rv8489b;      end
`else
`ifdef MODE_FORWARD
         assign jc52b77 = 1'b0;         assign ir95bbb = 1'b0;
`else
         assign jc52b77 = 1'b1;         assign ir95bbb = 1'b1;
`endif
`endif
`ifdef SFACT_PORT_READ
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ri9c793 <= {{`NUM_STAGES{2'b00}}};            lf137ce  <= {{`NUM_STAGES{2'b00}}};         end else begin            if(sfactset) ri9c793 <= sfact;            if(ibstart) begin               if(sfactset) lf137ce <= sfact;               else         lf137ce <= ri9c793 ;            end         end      end
`else
`endif
      assign qi2eb1c   = nga7d44>=ne5dba1 && kq5394e>=db288fc;
            always @(posedge clk or negedge rstn)      begin         if(!rstn) vx813b2 <= gb5451b;         else      vx813b2 <= ph9d96;      end
`ifdef BIT_REVERSE
      always @*      begin         case(vx813b2)            gb5451b     :  if(ibstart)             ph9d96 <= jea28dd;                        else                    ph9d96 <= gb5451b;            jea28dd    :  if(kq5394e>=db288fc)        ph9d96 <= pu146eb;                        else                    ph9d96 <= jea28dd;            pu146eb    :  if(kq5394e>=db288fc)        ph9d96 <= coa375b;                        else                    ph9d96 <= pu146eb;            coa375b     :  if(al65d63[`WR_LATENCY-1]) ph9d96 <= hq1bad8;                        else                    ph9d96 <= coa375b;            hq1bad8     :  if(qi2eb1c)                           if(ibstart)          ph9d96 <= jea28dd;                           else                 ph9d96 <= gb5451b;                        else                    ph9d96 <= hq1bad8;            default  :  ph9d96 <= gb5451b;         endcase      end
`else
      always @*      begin         case(vx813b2)            gb5451b     :  if(ibstart)             ph9d96 <= jea28dd;                        else                    ph9d96 <= gb5451b;            jea28dd    :  if(kq5394e>=db288fc)        ph9d96 <= pu146eb;                        else                    ph9d96 <= jea28dd;            pu146eb    :  if(kq5394e>=db288fc)        ph9d96 <= coa375b;                        else                    ph9d96 <= pu146eb;            coa375b     :  if(al65d63[`WR_LATENCY-1]) ph9d96 <= hq1bad8;                        else                    ph9d96 <= coa375b;            hq1bad8     :  if(qi2eb1c)            ph9d96 <= ym1f53c;                        else                    ph9d96 <= hq1bad8;            ym1f53c  :  if(tjb0a23>=db288fc)        ph9d96 <= wwfa9e0;                        else                    ph9d96 <= ym1f53c;            wwfa9e0  :  if(tjb0a23>=db288fc)                           if(ibstart)          ph9d96 <= jea28dd;                           else                 ph9d96 <= gb5451b;                        else                    ph9d96 <= wwfa9e0;            default  :  ph9d96 <= gb5451b;         endcase      end
`endif
      assign yx758e1 = (vx813b2==jea28dd)||(vx813b2==pu146eb)||(vx813b2==hq1bad8);
`ifdef BIT_REVERSE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                          nrf9dba <= 1'b0;         else if(db1c34b && tjb0a23>=db288fc) nrf9dba <= 1'b1;         else if(!db1c34b)                nrf9dba <= 1'b0;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                        db1c34b <= 1'b0;         else if(qi2eb1c)                db1c34b <= 1'b1;         else if(tjb0a23>=db288fc && nrf9dba) db1c34b <= 1'b0;      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                                 db1c34b <= 1'b0;         else if(qi2eb1c)                         db1c34b <= 1'b1;         else if(tjb0a23>=db288fc && vx813b2==wwfa9e0) db1c34b <= 1'b0;      end
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                                 rg63869 <= 1'b0;         else if(vx813b2==pu146eb && kq5394e>=db288fc)   rg63869 <= 1'b1;         else if(uv54fa8>=ne5dba1 && tjb0a23>=db288fc) rg63869 <= 1'b0;      end
      assign xj50aed = vx813b2==jea28dd || vx813b2==pu146eb;
      assign mgac70d = rg63869 || db1c34b;
      assign mt8576e = db1c34b;
      always @(posedge clk or negedge rstn)      begin         if(!rstn) for(en75165=0;en75165<`WR_LATENCY;en75165=en75165+1) al65d63[en75165] <= 1'b0;         else begin            al65d63[0] <= kq5394e>=db288fc;            for(en75165=1;en75165<`WR_LATENCY;en75165=en75165+1) al65d63[en75165] <=  al65d63[en75165-1];         end      end
      assign wj5142b = vx813b2==hq1bad8;      assign ir8a15d = rg63869;
      always @(posedge clk or negedge rstn)      begin         if(!rstn)      tjb0a23 <= {`LOG2_NBY2{1'b0}};         else if(mgac70d) tjb0a23 <= tjb0a23 + sw2bb74;         else           tjb0a23 <= {`LOG2_NBY2{1'b0}};      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)      kq5394e <= {`LOG2_NBY2{1'b0}};         else if(yx758e1) kq5394e <= kq5394e + sw2bb74;         else           kq5394e <= {`LOG2_NBY2{1'b0}};      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn)                  uv54fa8 <= {`STAGE_WIDTH{1'b0}};         else if(vx813b2==hq1bad8)            if(tjb0a23>=db288fc)               if(uv54fa8>=ne5dba1) uv54fa8 <= {`STAGE_WIDTH{1'b0}};               else                 uv54fa8 <= uv54fa8 + 1'b1;            else               uv54fa8 <= uv54fa8;         else                       uv54fa8 <= {`STAGE_WIDTH{1'b0}};      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                  nga7d44 <= {`STAGE_WIDTH{1'b0}};         else if(vx813b2==hq1bad8)            if(kq5394e>=db288fc)               if(nga7d44>=ne5dba1) nga7d44 <= {`STAGE_WIDTH{1'b0}};               else                 nga7d44 <= nga7d44 + 1'b1;            else               nga7d44 <= nga7d44;         else                       nga7d44 <= {`STAGE_WIDTH{1'b0}};      end
      
`ifdef BIT_REVERSE
`ifdef DYNAMIC_POINTS
         always @(posedge clk or negedge rstn)         begin            if(!rstn)        rfib <= 1'b1;            else if(ibstart) rfib <= 1'b0;            else if((!uv447e6[ri2a8a3-2] && uv447e6[ri2a8a3-3] && (ne5dba1==ym1a686)) ||                    (uv447e6[ri2a8a3-1] && !uv447e6[ri2a8a3-2] && vx813b2!=jea28dd && vx813b2!=pu146eb))               rfib <= 1'b1;         end
`else
         always @(posedge clk or negedge rstn)         begin            if(!rstn)        rfib <= 1'b1;            else if(ibstart) rfib <= 1'b0;            else if((!uv447e6[ri2a8a3-2] && uv447e6[ri2a8a3-3]) ||                    (uv447e6[ri2a8a3-1] && !uv447e6[ri2a8a3-2] && vx813b2!=jea28dd && vx813b2!=pu146eb))               rfib <= 1'b1;         end
`endif
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                                 rfib <= 1'b1;         else if(ibstart)                          rfib <= 1'b0;         else if(vx813b2==wwfa9e0 && tjb0a23>=db288fc) rfib <= 1'b1;      end
`endif
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            dz5f51c     <= 1'b0;            rg697d4 <= 1'b0;            gb4bea3 <= 1'b0;            vka88c0     <= 1'b0;            ip44602     <= 1'b0;         end else begin            dz5f51c     <= vx813b2==hq1bad8;            rg697d4 <= vx813b2==jea28dd || dz5f51c;            gb4bea3 <= vx813b2==pu146eb || dz5f51c;            vka88c0     <= rg697d4;            ip44602     <= gb4bea3;         end      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            kqfa8e6 <= {(`WR_LATENCY+1){1'b0}};            swa3981 <= {(`WR_LATENCY+2){1'b0}};         end else begin            kqfa8e6 <= {kqfa8e6[`WR_LATENCY-1:0],rg63869};            swa3981 <= {swa3981[`WR_LATENCY:0],uv54fa8>=ne5dba1};         end      end      always @(posedge clk or negedge rstn)      begin         if(!rstn)                       pf742a7 <= 1'b0;         else if(kqfa8e6[`WR_LATENCY]) pf742a7 <= ~pf742a7;         else                            pf742a7 <= 1'b0;      end
`ifdef TRUNCATE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                         uka9d85 <= 1'b0;         else if(kqfa8e6[`WR_LATENCY-4]) uka9d85 <= ~uka9d85;         else                              uka9d85 <= 1'b0;      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)                         uka9d85 <= 1'b0;         else if(kqfa8e6[`WR_LATENCY-5]) uka9d85 <= ~uka9d85;         else                              uka9d85 <= 1'b0;      end
`endif
      assign qva153e = swa3981[`WR_LATENCY+1];
            always @(posedge clk or negedge rstn)      begin         if(!rstn) uk3ea23 <= 1'b0;         else      uk3ea23 <= xj50aed;      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) uv447e6 <= {ri2a8a3{1'b0}};         else      uv447e6 <= {uv447e6[ri2a8a3-2:0],db1c34b};      end
      assign vica285 = uv447e6[3];
`ifdef TRUNCATE
      assign outvalid = uv447e6[7];      assign uvd9450   = uv447e6[6];
`else
      assign outvalid = uv447e6[8];      assign uvd9450 = uv447e6[7];
`endif
      
`ifdef OUTVALID_SEL
`ifdef TRUNCATE
           assign ng14954 = uv447e6[5];
`else
           assign ng14954 = uv447e6[6];
`endif
`endif
   
      
`ifdef TRUNCATE
      always @(posedge clk or negedge rstn)      begin         if(!rstn) obstart <= 1'b0;         else      obstart <= !uv447e6[7] && uv447e6[6];      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) obstart <= 1'b0;         else      obstart <= !uv447e6[8] && uv447e6[7];      end
`endif
            always @(posedge clk or negedge rstn)      begin         if(!rstn) je30276 <= 8'h01;         else begin            if(mt8576e && tjb0a23>=db288fc) je30276[0] <= 1'b0;            else if(!mt8576e)           je30276[0] <= 1'b1;            je30276[7:1] <= {je30276[6:1],je30276[0]};         end      end
`ifdef TRUNCATE
      assign gof5118 = je30276[6];
`else
      assign gof5118 = je30276[7];
`endif
            always @(posedge clk or negedge rstn)      begin         if(!rstn) ibend <= 1'b0;         else      ibend <= (kq5394e==(`NUM_POINTS/2 - {sw2bb74,2'b00}))&& (vx813b2==pu146eb);      end
            assign al4ec28 = rg63869;      assign fa76144  = uv447e6[2];      assign qi1f9a5 = uv447e6[3];      assign oh23014 = ibend;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
      
`ifdef SFACT_PORT_READ
`ifdef NUM_POINTS_64
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];               endcase            end
`endif
`ifdef NUM_POINTS_128
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];               endcase            end
`endif
`ifdef NUM_POINTS_256
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];               endcase            end
`endif
`ifdef NUM_POINTS_512
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];               endcase            end
`endif
`ifdef NUM_POINTS_1024
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];                  9  :  cz709f8 <= lf137ce[`SFACT_WIDTH-19:`SFACT_WIDTH-20];               endcase            end
`endif
`ifdef NUM_POINTS_2048
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];                  9  :  cz709f8 <= lf137ce[`SFACT_WIDTH-19:`SFACT_WIDTH-20];                  10 :  cz709f8 <= lf137ce[`SFACT_WIDTH-21:`SFACT_WIDTH-22];               endcase            end
`endif
`ifdef NUM_POINTS_4096
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];                  9  :  cz709f8 <= lf137ce[`SFACT_WIDTH-19:`SFACT_WIDTH-20];                  10 :  cz709f8 <= lf137ce[`SFACT_WIDTH-21:`SFACT_WIDTH-22];                  11 :  cz709f8 <= lf137ce[`SFACT_WIDTH-23:`SFACT_WIDTH-24];               endcase            end
`endif
`ifdef NUM_POINTS_8192
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];                  9  :  cz709f8 <= lf137ce[`SFACT_WIDTH-19:`SFACT_WIDTH-20];                  10 :  cz709f8 <= lf137ce[`SFACT_WIDTH-21:`SFACT_WIDTH-22];                  11 :  cz709f8 <= lf137ce[`SFACT_WIDTH-23:`SFACT_WIDTH-24];                  12 :  cz709f8 <= lf137ce[`SFACT_WIDTH-25:`SFACT_WIDTH-26];               endcase            end
`endif
`ifdef NUM_POINTS_16384
            always @(posedge clk or negedge rstn)            begin               if(!rstn) cz709f8 <= 2'b00;               else case(uv54fa8)                  0  :  cz709f8 <= lf137ce[`SFACT_WIDTH-1:`SFACT_WIDTH-2];                  1  :  cz709f8 <= lf137ce[`SFACT_WIDTH-3:`SFACT_WIDTH-4];                  2  :  cz709f8 <= lf137ce[`SFACT_WIDTH-5:`SFACT_WIDTH-6];                  3  :  cz709f8 <= lf137ce[`SFACT_WIDTH-7:`SFACT_WIDTH-8];                  4  :  cz709f8 <= lf137ce[`SFACT_WIDTH-9:`SFACT_WIDTH-10];                  5  :  cz709f8 <= lf137ce[`SFACT_WIDTH-11:`SFACT_WIDTH-12];                  6  :  cz709f8 <= lf137ce[`SFACT_WIDTH-13:`SFACT_WIDTH-14];                  7  :  cz709f8 <= lf137ce[`SFACT_WIDTH-15:`SFACT_WIDTH-16];                  8  :  cz709f8 <= lf137ce[`SFACT_WIDTH-17:`SFACT_WIDTH-18];                  9  :  cz709f8 <= lf137ce[`SFACT_WIDTH-19:`SFACT_WIDTH-20];                  10 :  cz709f8 <= lf137ce[`SFACT_WIDTH-21:`SFACT_WIDTH-22];                  11 :  cz709f8 <= lf137ce[`SFACT_WIDTH-23:`SFACT_WIDTH-24];                  12 :  cz709f8 <= lf137ce[`SFACT_WIDTH-25:`SFACT_WIDTH-26];                  13 :  cz709f8 <= lf137ce[`SFACT_WIDTH-27:`SFACT_WIDTH-28];               endcase            end
`endif
         always @(posedge clk or negedge rstn)         begin            if(!rstn)               for(en75165=0;en75165<`WR_LATENCY;en75165=en75165+1) bab84f6[en75165] <= 2'b00;            else begin               bab84f6[0] <= cz709f8;               for(en75165=1;en75165<`WR_LATENCY;en75165=en75165+1) bab84f6[en75165] <= bab84f6[en75165-1];            end         end
`ifdef TRUNCATE
         always @(posedge clk or negedge rstn)         begin            if(!rstn)          aaacedc <= 2'b00;            else if(uv447e6[3]) aaacedc <= 2'b00;            else               aaacedc <= bab84f6[`WR_LATENCY-3];         end
`else
         always @(posedge clk or negedge rstn)         begin            if(!rstn)          aaacedc <= 2'b00;            else if(uv447e6[3]) aaacedc <= 2'b00;            else               aaacedc <= bab84f6[`WR_LATENCY-4];         end
`endif
`endif
`ifdef SFACT_UNSCALE
`endif
`ifdef SFACT_RS111
         always @(posedge clk or negedge rstn)         begin            if(!rstn)          aaacedc <= 2'b00;            else if(qi1f9a5) aaacedc <= 2'b00;            else               aaacedc <= 2'b01;         end
`endif
`ifdef SFACT_RS211
         always @(posedge clk or negedge rstn)         begin            if(!rstn)               for(en75165=0;en75165<`WR_LATENCY;en75165=en75165+1) pff65ff[en75165] <= 1'b0;            else begin               pff65ff[0] <= uv54fa8=={`STAGE_WIDTH{1'b0}};               for(en75165=1;en75165<`WR_LATENCY;en75165=en75165+1) pff65ff[en75165] <= pff65ff[en75165-1];            end         end
`ifdef TRUNCATE
            always @(posedge clk or negedge rstn)            begin               if(!rstn)                       aaacedc <= 2'b00;               else if(qi1f9a5)              aaacedc <= 2'b00;               else if(pff65ff[`WR_LATENCY-2]) aaacedc <= 2'b10;               else                            aaacedc <= 2'b01;            end
`else
            always @(posedge clk or negedge rstn)            begin               if(!rstn)                       aaacedc <= 2'b00;               else if(qi1f9a5)              aaacedc <= 2'b00;               else if(pff65ff[`WR_LATENCY-3]) aaacedc <= 2'b10;               else                            aaacedc <= 2'b01;            end
`endif
`endif
                  always @(posedge clk or negedge rstn)         begin            if(!rstn)                               by76eb8 <= 1'b0;            else if(vx813b2==pu146eb && kq5394e>=db288fc) by76eb8 <= 1'b0;            else                                    by76eb8 <= by76eb8 || dmfb548;         end
`ifdef TRUNCATE
         always @(posedge clk or negedge rstn)         begin            if(!rstn)          except <= 1'b0;            else if(uv447e6[6]) except <= by76eb8;            else               except <= 1'b0;         end
`else
         always @(posedge clk or negedge rstn)         begin            if(!rstn)          except <= 1'b0;            else if(uv447e6[7]) except <= by76eb8;            else               except <= 1'b0;         end
`endif
`endif
`endif
   endmodule                                                                                                   
`timescale 1 ns / 100 ps
module epd4c0_FFTC2048 (
               rstn,             
               clk,              
               aa98120,              
   
   
           `ifdef OUTVALID_SEL
               ng14954,
           `endif
   
               rv2dca9,            
               dz6e54e,            
               su72a76,            
               oh953b0,            
   
               dore,             
               doim              
            );
input                   rstn;
input                   clk;
input                   aa98120;
`ifdef OUTVALID_SEL
input                   ng14954;
`endif
input [`DATA_WIDTH-1:0] rv2dca9;
input [`DATA_WIDTH-1:0] dz6e54e;
input [`DATA_WIDTH-1:0] su72a76;
input [`DATA_WIDTH-1:0] oh953b0;
output[`DATA_WIDTH-1:0] dore;
output[`DATA_WIDTH-1:0] doim;
reg [`DATA_WIDTH-1:0]   dore;
reg [`DATA_WIDTH-1:0]   doim;
`ifdef OUTVALID_SEL
`else
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef OUTVALID_SEL
`else
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef OUTVALID_SEL
`else
`endif
         
`ifdef OUTVALID_SEL
`endif
            
`ifdef OUTVALID_SEL
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            dore <= {`DATA_WIDTH{1'b0}};            doim <= {`DATA_WIDTH{1'b0}};         end else begin             case({ng14954,aa98120})                 2'b10: begin                           dore <= su72a76;                           doim <= oh953b0;                        end                 2'b11: begin                           dore <= rv2dca9;                           doim <= dz6e54e;                        end                 default: begin                           dore <= {`DATA_WIDTH{1'b0}};                           doim <= {`DATA_WIDTH{1'b0}};                        end             endcase         end      end
`else
         always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            dore <= {`DATA_WIDTH{1'b0}};            doim <= {`DATA_WIDTH{1'b0}};         end else if(aa98120) begin            dore <= rv2dca9;            doim <= dz6e54e;         end else begin            dore <= su72a76;            doim <= oh953b0;         end      end
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module sj232d3_FFTC2048 (
               rstn,                
               clk,                 
               uk3ea23,                
               end39ce,           
               tw9ce75,           
               rv2dca9,               
               dz6e54e,               
               su72a76,               
               oh953b0,               
               pf742a7,               
               qva153e,               
               ks34a7f,               
               hda53f9,               
               an29fcf,               
               xj4fe7c                
               );
input                      rstn;
input                      clk;
input                      uk3ea23;
input [`DATA_WIDTH-1:0]    end39ce;
input [`DATA_WIDTH-1:0]    tw9ce75;
input [`DATA_WIDTH-1:0]    rv2dca9;
input [`DATA_WIDTH-1:0]    dz6e54e;
input [`DATA_WIDTH-1:0]    su72a76;
input [`DATA_WIDTH-1:0]    oh953b0;
input                      pf742a7;
input                      qva153e;
output[`DATA_WIDTH-1:0]    ks34a7f;
output[`DATA_WIDTH-1:0]    hda53f9;
output[`DATA_WIDTH-1:0]    an29fcf;
output[`DATA_WIDTH-1:0]    xj4fe7c;
reg [`DATA_WIDTH-1:0]      ks34a7f;
reg [`DATA_WIDTH-1:0]      hda53f9;
reg [`DATA_WIDTH-1:0]      an29fcf;
reg [`DATA_WIDTH-1:0]      xj4fe7c;
reg [`DATA_WIDTH-1:0]      ohd391;
reg [`DATA_WIDTH-1:0]      ne69c8c;
reg [`DATA_WIDTH-1:0]      wj4e462;
reg [`DATA_WIDTH-1:0]      cm72315;
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ohd391 <= {(`DATA_WIDTH){1'b0}};            ne69c8c <= {(`DATA_WIDTH){1'b0}};            wj4e462 <= {(`DATA_WIDTH){1'b0}};            cm72315 <= {(`DATA_WIDTH){1'b0}};         end else if(pf742a7 && !qva153e) begin            ohd391 <= su72a76;            ne69c8c <= oh953b0;         end else begin            ohd391 <= rv2dca9;            ne69c8c <= dz6e54e;            wj4e462 <= su72a76;            cm72315 <= oh953b0;         end      end
            always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ks34a7f <= {(`DATA_WIDTH){1'b0}};            hda53f9 <= {(`DATA_WIDTH){1'b0}};            an29fcf <= {(`DATA_WIDTH){1'b0}};            xj4fe7c <= {(`DATA_WIDTH){1'b0}};         end else if(uk3ea23) begin            ks34a7f <= end39ce;            hda53f9 <= tw9ce75;            an29fcf <= end39ce;            xj4fe7c <= tw9ce75;         end else if(qva153e) begin            ks34a7f <= ohd391;            hda53f9 <= ne69c8c;            an29fcf <= wj4e462;            xj4fe7c <= cm72315;         end else if(pf742a7) begin            ks34a7f <= ohd391;            hda53f9 <= ne69c8c;            an29fcf <= rv2dca9;            xj4fe7c <= dz6e54e;         end else begin            ks34a7f <= wj4e462;            hda53f9 <= cm72315;            an29fcf <= ohd391;            xj4fe7c <= ne69c8c;         end      end
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module rtf9aaf_FFTC2048 (
               rstn,                
               clk,                 
               vica285,            
               cz709f8,              
               rv2dca9,               
               dz6e54e,               
               su72a76,               
               oh953b0,               
               go7788d,
               ukbc468,
               ipe2340,
               do11a04,
            `ifdef BFPU_PRESENT
            `else
            `ifdef SFACT_UNSCALE
            `else
               except,              
            `endif
            `endif
               ks34a7f,               
               hda53f9,               
               an29fcf,               
               xj4fe7c                
            );
input                      rstn;
input                      clk;
input                      vica285;
input [1:0]                cz709f8;
input [`DATA_WIDTH+1:0]    rv2dca9;
input [`DATA_WIDTH+1:0]    dz6e54e;
input [`DATA_WIDTH+1:0]    su72a76;
input [`DATA_WIDTH+1:0]    oh953b0;
input [`DATA_WIDTH-1:0]    go7788d;
input [`DATA_WIDTH-1:0]    ukbc468;
input [`DATA_WIDTH-1:0]    ipe2340;
input [`DATA_WIDTH-1:0]    do11a04;
output[`DATA_WIDTH-1:0]    ks34a7f;
output[`DATA_WIDTH-1:0]    hda53f9;
output[`DATA_WIDTH-1:0]    an29fcf;
output[`DATA_WIDTH-1:0]    xj4fe7c;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
output                     except;
reg                        except;
wire                       ldfcc78;
wire                       the63c7;
wire                       mg31e3e;
wire                       wl8f1f1;
`endif
`endif
wire[`DATA_WIDTH+1:0]      ksf3af;
wire[`DATA_WIDTH+1:0]      lq79d79;
wire[`DATA_WIDTH+1:0]      qgcebcb;
wire[`DATA_WIDTH+1:0]      en75e58;
wire[1:0]                  cz709f8;
reg                        fa7962e;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) fa7962e <= 1'b0;         else      fa7962e <= vica285;      end
      assign ksf3af = fa7962e ? {{2{go7788d[`DATA_WIDTH-1]}},go7788d} : rv2dca9;      assign lq79d79 = fa7962e ? {{2{ukbc468[`DATA_WIDTH-1]}},ukbc468} : dz6e54e;      assign qgcebcb = fa7962e ? {{2{ipe2340[`DATA_WIDTH-1]}},ipe2340} : su72a76;      assign en75e58 = fa7962e ? {{2{do11a04[`DATA_WIDTH-1]}},do11a04} : oh953b0;
      vxb030e_FFTC2048 nt81876 (               .clk        (clk         ),               .rstn       (rstn        ),               .din        (ksf3af      ),               .cz709f8      (cz709f8       ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
               .except     (ldfcc78  ),
`endif
`endif
               .dout       (ks34a7f       )              ) ;
      vxb030e_FFTC2048 hbd8391 (               .clk        (clk         ),               .rstn       (rstn        ),               .din        (lq79d79      ),               .cz709f8      (cz709f8       ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
               .except     (the63c7  ),
`endif
`endif
               .dout       (hda53f9       )              ) ;
      vxb030e_FFTC2048 ld409a8 (               .clk        (clk         ),               .rstn       (rstn        ),               .din        (qgcebcb      ),               .cz709f8      (cz709f8       ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
               .except     (mg31e3e  ),
`endif
`endif
               .dout       (an29fcf       )              ) ;
      vxb030e_FFTC2048 nrc243e (               .clk        (clk         ),               .rstn       (rstn        ),               .din        (en75e58      ),               .cz709f8      (cz709f8       ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
               .except     (wl8f1f1  ),
`endif
`endif
               .dout       (xj4fe7c       )              ) ;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) except <= 1'b0;         else      except <= ldfcc78 | the63c7 | mg31e3e | wl8f1f1;      end
`endif
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module vxb030e_FFTC2048 (
            clk,                  
            rstn,                 
            din,                  
            cz709f8,                
         `ifdef BFPU_PRESENT
         `else
         `ifdef SFACT_UNSCALE
         `else
            except,               
         `endif
         `endif
            dout                  
          ) ;
input                      clk;
input                      rstn;
input [`DATA_WIDTH+1:0]    din;
input [1:0]                cz709f8;
output [`DATA_WIDTH-1:0]   dout;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
output                     except;
`endif
`endif
reg [`DATA_WIDTH-1:0]      dout;
wire                       ne57a3b;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
reg                        except;
`endif
`endif
`ifdef TRUNCATE
reg [`DATA_WIDTH-1:0] sue069f;
`else
reg [`DATA_WIDTH-1:0]   lf34f9;
reg                     shfd9a1;
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef TRUNCATE
`else
`endif
            
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
                  assign ne57a3b = din[`DATA_WIDTH+1] ;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            except <= 1'b0;         else case(cz709f8)            2'b00   : except <= (|din[`DATA_WIDTH+1:`DATA_WIDTH-1])&(!(&din[`DATA_WIDTH+1:`DATA_WIDTH-1]));            2'b01   : except <= (|din[`DATA_WIDTH+1:`DATA_WIDTH])&(!(&din[`DATA_WIDTH+1:`DATA_WIDTH]));            default : except <= 1'b0;         endcase      end
`endif
`endif
`ifdef TRUNCATE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            dout <= {`DATA_WIDTH{1'b0}};         else case(cz709f8)            2'b00   : dout <= {ne57a3b,din[`DATA_WIDTH-2:0]};            2'b01   : dout <= {ne57a3b,din[`DATA_WIDTH-1:1]};            2'b10   : dout <= {ne57a3b,din[`DATA_WIDTH:2]};            default : dout <= {ne57a3b,din[`DATA_WIDTH-2:0]};         endcase      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            lf34f9 <= {`DATA_WIDTH{1'b0}};            shfd9a1    <= 1'b0;         end else case(cz709f8)            2'b00 :  begin                        lf34f9 <= {ne57a3b,din[`DATA_WIDTH-2:0]};                        shfd9a1    <= 1'b0;                     end            2'b01 :  begin                        lf34f9 <= {ne57a3b,din[`DATA_WIDTH-1:1]};                        shfd9a1 <= ne57a3b ? 1'b0 : din[0];                     end            2'b10 :  begin                        lf34f9 <= {ne57a3b,din[`DATA_WIDTH:2]};                        shfd9a1 <= ne57a3b ? (&din[1:0]) : din[1];                     end            default : begin                        lf34f9 <= {ne57a3b,din[`DATA_WIDTH-2:0]};                        shfd9a1    <= 1'b0;                      end         endcase      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) dout <= {`DATA_WIDTH{1'b0}};         else      dout <= lf34f9 + shfd9a1;      end
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module yx4b493_FFTC2048 (
                  rstn,             
                  clk,              
                  tjb0a23,             
                  uv54fa8,           
               `ifdef TMEM_ALL
               `else
                  qi9dd83,        
                  lqeec18,           
               `endif
                  jc760c3            
               ) ;
input                      rstn;
input                      clk;
input [`LOG2_NBY2-1:0]     tjb0a23;
input [`STAGE_WIDTH-1:0]   uv54fa8;
`ifdef TMEM_ALL
output[`LOG2_NBY2-1:0]     jc760c3;
`else
output[1:0]                qi9dd83;
output[`LOG2_NBY4-1:0]     lqeec18;
output[`LOG2_NBY4-1:0]     jc760c3;
`endif
`ifdef TMEM_ALL
reg [`LOG2_NBY2-1:0]       jc760c3;
`else
reg [`LOG2_NBY4-1:0]       lqeec18;
reg [1:0]                  qi9dd83;
reg [1:0]                  yxc6172[0:1];
reg [`LOG2_NBY4-1:0]       jc760c3;
`endif
reg [`LOG2_NBY2-1:0]       ux85cab;
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TMEM_ALL
reg [`LOG2_NBY2-1:0] ie2e55d;
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
      
`ifdef NUM_POINTS_64
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_128
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_256
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_512
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_1024
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-8],{(`LOG2_NBY2-8){1'b0}}};            9  :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_2048
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-8],{(`LOG2_NBY2-8){1'b0}}};            9  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-9],{(`LOG2_NBY2-9){1'b0}}};            10 :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_4096
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-8],{(`LOG2_NBY2-8){1'b0}}};            9  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-9],{(`LOG2_NBY2-9){1'b0}}};            10 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-10],{(`LOG2_NBY2-10){1'b0}}};            11 :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_8192
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-8],{(`LOG2_NBY2-8){1'b0}}};            9  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-9],{(`LOG2_NBY2-9){1'b0}}};            10 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-10],{(`LOG2_NBY2-10){1'b0}}};            11 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-11],{(`LOG2_NBY2-11){1'b0}}};            12 :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef NUM_POINTS_16384
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ux85cab <= {`LOG2_NBY2{1'b0}};         else case(uv54fa8)            0  :  ux85cab <= {`LOG2_NBY2{1'b0}};            1  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1],{(`LOG2_NBY2-1){1'b0}}};            2  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-2],{(`LOG2_NBY2-2){1'b0}}};            3  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-3],{(`LOG2_NBY2-3){1'b0}}};            4  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-4],{(`LOG2_NBY2-4){1'b0}}};            5  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-5],{(`LOG2_NBY2-5){1'b0}}};            6  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-6],{(`LOG2_NBY2-6){1'b0}}};            7  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-7],{(`LOG2_NBY2-7){1'b0}}};            8  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-8],{(`LOG2_NBY2-8){1'b0}}};            9  :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-9],{(`LOG2_NBY2-9){1'b0}}};            10 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-10],{(`LOG2_NBY2-10){1'b0}}};            11 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-11],{(`LOG2_NBY2-11){1'b0}}};            12 :  ux85cab <= {tjb0a23[`LOG2_NBY2-1:`LOG2_NBY2-12],{(`LOG2_NBY2-12){1'b0}}};            13 :  ux85cab <= tjb0a23;            default : ux85cab <= tjb0a23;         endcase      end
`endif
`ifdef TMEM_ALL
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ie2e55d <= {`LOG2_NBY2{1'b0}};            jc760c3     <= {`LOG2_NBY2{1'b0}};         end else begin            ie2e55d <= ux85cab;            jc760c3     <= ie2e55d;         end      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            jc760c3           <= {`LOG2_NBY4{1'b0}};            lqeec18           <= {`LOG2_NBY4{1'b0}};            yxc6172[0] <= 2'b00;         end else if(ux85cab==0) begin            jc760c3           <= {`LOG2_NBY4{1'b0}};            lqeec18           <= {`LOG2_NBY4{1'b0}};            yxc6172[0] <= 2'b00;         end else if(ux85cab==`NUM_POINTS/4) begin            jc760c3           <= {`LOG2_NBY4{1'b0}};            lqeec18           <= {`LOG2_NBY4{1'b0}};            yxc6172[0] <= 2'b01;         end else if(ux85cab < `NUM_POINTS/4) begin            jc760c3           <= ux85cab;            lqeec18           <= `NUM_POINTS/4 - ux85cab;            yxc6172[0] <= 2'b10;         end else begin            jc760c3           <= `NUM_POINTS/4 - ux85cab;            lqeec18           <= ux85cab - `NUM_POINTS/4;            yxc6172[0] <= 2'b11;         end      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            qi9dd83        <= 2'b00;            yxc6172[1] <= 2'b00;         end else begin            yxc6172[1] <= yxc6172[0];            qi9dd83        <= yxc6172[1];         end      end
`endif
   endmodule                                                                                             
`timescale 1 ns / 100 ps
module dmfb478_FFTC2048 (
               clk,              
               rstn,             
               jc760c3,           
            `ifdef TMEM_ALL
            `else
               lqeec18,           
               qi9dd83,        
            `endif
               aa1a145             
               );
input                      clk;
input                      rstn;
`ifdef TMEM_ALL
input [`LOG2_NBY2-1:0]     jc760c3;
`else
input [`LOG2_NBY4-1:0]     lqeec18;
input [1:0]                qi9dd83;
input [`LOG2_NBY4-1:0]     jc760c3;
`endif
output[`TWID_WIDTH2-1:0]   aa1a145;
`ifdef USE_DIST_ROM
wire[`TWID_WIDTH2-1:0]        eca6dd2;
reg [`TWID_WIDTH2-1:0]        aa1a145;
`else
`ifdef TMEM_ALL
`else
wire [`TWID_WIDTH-1:0]    mt293f0;
wire [`TWID_WIDTH-1:0]    jp4fc29;
reg  [`TWID_WIDTH-1:0]    vvd231f;
reg  [`TWID_WIDTH-1:0]    xl918fe;
`endif
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef USE_DIST_ROM
`else
`ifdef TMEM_ALL
`else
`endif
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef USE_DIST_ROM
`else
`ifdef TMEM_ALL
`else
`endif
`endif
      
`ifdef TMEM_ALL
`else
`endif
      
`ifdef USE_DIST_ROM
      defparam ls8c7f6.pmi_addr_depth       = (`NUM_POINTS/2);      defparam ls8c7f6.pmi_addr_width       = (`LOG2_N-1);      defparam ls8c7f6.pmi_data_width       = `TWID_WIDTH2;      defparam ls8c7f6.pmi_regmode          = "reg";      defparam ls8c7f6.pmi_init_file        = "twidFFTC2048.mem";      defparam ls8c7f6.pmi_init_file_format = "binary";      defparam ls8c7f6.pmi_family           = `DEVICE_FAMILY;      defparam ls8c7f6.module_type          = "pmi_distributed_rom";      pmi_distributed_rom ls8c7f6 (                                 .Address    (jc760c3        ),                                 .OutClock   (clk           ),                                 .OutClockEn (1'b1          ),                                 .Reset      (1'b0          ),                                 .Q          (eca6dd2         )                              );
      always @(posedge clk or negedge rstn)      begin         if(!rstn) aa1a145 <= {`TWID_WIDTH2{1'b0}};         else      aa1a145 <= eca6dd2;      end
`else
`ifdef TMEM_ALL
         defparam suf55ba.pmi_addr_depth = (`NUM_POINTS/2);         defparam suf55ba.pmi_addr_width = (`LOG2_N-1);         defparam suf55ba.pmi_data_width = `TWID_WIDTH2;         defparam suf55ba.pmi_regmode = "reg";         defparam suf55ba.pmi_gsr = "disable";         defparam suf55ba.pmi_resetmode = "sync";         defparam suf55ba.pmi_init_file = "twidFFTC2048.mem";         defparam suf55ba.pmi_init_file_format = "binary";         defparam suf55ba.pmi_family = `DEVICE_FAMILY;         defparam suf55ba.module_type = "pmi_rom";         pmi_rom suf55ba (                           .Address       (jc760c3     ),                           .OutClock      (clk        ),                           .OutClockEn    (1'b1       ),                           .Reset         (1'b0       ),                           .Q             (aa1a145      )                        );
`else
         defparam zkf1fa0.pmi_addr_depth_a = `NBY4;         defparam zkf1fa0.pmi_addr_width_a = `LOG2_NBY4;         defparam zkf1fa0.pmi_data_width_a = `TWID_WIDTH;         defparam zkf1fa0.pmi_addr_depth_b = `NBY4;         defparam zkf1fa0.pmi_addr_width_b = `LOG2_NBY4;         defparam zkf1fa0.pmi_data_width_b = `TWID_WIDTH;         defparam zkf1fa0.pmi_regmode_a = "reg";         defparam zkf1fa0.pmi_regmode_b = "reg";         defparam zkf1fa0.pmi_gsr = "disable";         defparam zkf1fa0.pmi_resetmode = "sync";         defparam zkf1fa0.pmi_init_file = "twidFFTC2048.mem";         defparam zkf1fa0.pmi_init_file_format = "binary";         defparam zkf1fa0.pmi_write_mode_a = "normal";         defparam zkf1fa0.pmi_write_mode_b = "normal";         defparam zkf1fa0.pmi_family = `DEVICE_FAMILY;         defparam zkf1fa0.module_type = "pmi_ram_dp_true";         pmi_ram_dp_true zkf1fa0 (                           .DataInA    (           ),                           .DataInB    (           ),                           .AddressA   (jc760c3     ),                           .AddressB   (lqeec18     ),                           .ClockA     (clk        ),                           .ClockB     (clk        ),                           .ClockEnA   (1'b1       ),                           .ClockEnB   (1'b1       ),                           .WrA        (1'b0       ),                           .WrB        (1'b0       ),                           .ResetA     (1'b0       ),                           .ResetB     (1'b0       ),                           .QA         (mt293f0  ),                           .QB         (jp4fc29  )                        );
         always @(posedge clk or negedge rstn)         begin            if(!rstn) begin               vvd231f <= {`TWID_WIDTH{1'b0}};               xl918fe <= {`TWID_WIDTH{1'b0}};            end else begin               case(qi9dd83)                  2'b00 :  begin                              vvd231f <= mt293f0;                              xl918fe <= {`TWID_WIDTH{1'b0}};                           end                  2'b01 :  begin                              vvd231f <= {`TWID_WIDTH{1'b0}};                              xl918fe <= ~jp4fc29 + 1;                           end                  2'b10 :  begin                              vvd231f <= mt293f0;                              xl918fe <= ~jp4fc29 + 1;                           end                  2'b11 :  begin                              vvd231f <= ~mt293f0 + 1;                              xl918fe <= ~jp4fc29 + 1;                           end               endcase            end         end
         assign aa1a145 = {vvd231f,xl918fe};
`endif
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module ba2adc0_FFTC2048 (
                  rstn,                
                  clk,                 
                  ir8a15d,             
                  wj5142b,             
                  xj50aed,           
                  mt8576e,             
                  fn6e854,              
                  ne5dba1,
   
                  uv54fa8,              
               `ifdef BIT_REVERSE
                  an8511f,
               `endif
               `ifdef ADDRESS_OUT
                  oaddr,               
               `endif
                  thf9dcf,          
                  cmcee7f           
               );
input                      rstn;
input                      clk;
input [`STAGE_WIDTH-1:0]   uv54fa8;
input                      ir8a15d;
input                      wj5142b;
input                      xj50aed;
input                      mt8576e;
input [3:0]                fn6e854;
input [`STAGE_WIDTH-1:0]   ne5dba1;
`ifdef BIT_REVERSE
output[`LOG2_NBY2-1:0]     an8511f;
`endif
`ifdef ADDRESS_OUT
output[`LOG2_N-1:0]     oaddr;
`endif
output[`LOG2_NBY2-1:0]     thf9dcf;
output[`LOG2_NBY2-1:0]     cmcee7f;
reg [`LOG2_NBY2-1:0]       thf9dcf;
reg [`LOG2_NBY2-1:0]       cmcee7f;
reg                        xy8cd0d;
integer                    en75165;
reg                        ec3435b;
reg                        gda1ad8;
reg [`LOG2_NBY2-1:0]       ohd6c4;
reg [`LOG2_NBY2-1:0]       pf6b624;
reg [`LOG2_NBY2-1:0]       an8511f;
wire[`LOG2_NBY2-1:0]       hbd8934;
wire[`LOG2_NBY2-1:0]       qgc49a6;
reg [`STAGE_WIDTH-1:0]     co24d31;
reg   ir26988;
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
reg qi5137,ip75347;
reg [`LOG2_NBY2-1:0] aa31148[0:`WR_LATENCY-1];
`ifdef BIT_REVERSE
wire[`LOG2_NBY2-1:0] ym88a40;
`endif
reg   vv45201;
reg   oh2900e;
`ifdef BIT_REVERSE
`else
`endif
`ifdef ADDRESS_OUT
reg [`LOG2_N-1:0] ho48075[0:6];
reg [1:0]         ld403aa;
wire[`LOG2_N-1:0] ls1d56 = {ohd6c4[`LOG2_NBY2-1:1],2'b11};
wire[`LOG2_N-1:0] ykdbf27     = ~{1'b0,ohd6c4[`LOG2_NBY2-1:1],1'b1};
wire[`LOG2_N-1:0] kq566a7 = {`LOG2_N{ld403aa[1]}};
wire[`LOG2_N-1:0] gd9a9c1 = {1'b0,cmcee7f};
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef BIT_REVERSE
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef ADDRESS_OUT
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef BIT_REVERSE
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef ADDRESS_OUT
`ifdef TRUNCATE
`else
`endif
`endif
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) co24d31 <= {`STAGE_WIDTH{1'b0}};         else      co24d31 <= uv54fa8;      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ir26988 <= 1'b0;            xy8cd0d     <= 1'b0;         end else begin            ir26988 <= xj50aed;            xy8cd0d     <= ir26988;         end      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            ec3435b <= 1'b0;            gda1ad8 <= 1'b0;         end else begin            ec3435b <= wj5142b || xj50aed;            gda1ad8 <= ir8a15d || mt8576e;         end      end
`ifdef NUM_POINTS_64
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else      ohd6c4 <= `NUM_POINTS/2-2;      end
`endif
`ifdef NUM_POINTS_128
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ohd6c4 <= `NUM_POINTS/2-1;         else if(ne5dba1==5) ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};         else                 ohd6c4 <= `NUM_POINTS/2-2;      end
`endif
`ifdef NUM_POINTS_256
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_512
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_1024
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            8  :  ohd6c4 <= {{(`LOG2_NBY2-8){1'b0}},{7{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_2048
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            8  :  ohd6c4 <= {{(`LOG2_NBY2-8){1'b0}},{7{1'b1}},1'b0};            9  :  ohd6c4 <= {{(`LOG2_NBY2-9){1'b0}},{8{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_4096
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            8  :  ohd6c4 <= {{(`LOG2_NBY2-8){1'b0}},{7{1'b1}},1'b0};            9  :  ohd6c4 <= {{(`LOG2_NBY2-9){1'b0}},{8{1'b1}},1'b0};            10 :  ohd6c4 <= {{(`LOG2_NBY2-10){1'b0}},{9{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_8192
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            8  :  ohd6c4 <= {{(`LOG2_NBY2-8){1'b0}},{7{1'b1}},1'b0};            9  :  ohd6c4 <= {{(`LOG2_NBY2-9){1'b0}},{8{1'b1}},1'b0};            10 :  ohd6c4 <= {{(`LOG2_NBY2-10){1'b0}},{9{1'b1}},1'b0};            11 :  ohd6c4 <= {{(`LOG2_NBY2-11){1'b0}},{10{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
`ifdef NUM_POINTS_16384
      always @(posedge clk or negedge rstn)      begin         if(!rstn) ohd6c4 <= `NUM_POINTS/2-1;         else case(ne5dba1)            5  :  ohd6c4 <= {{(`LOG2_NBY2-5){1'b0}},{4{1'b1}},1'b0};            6  :  ohd6c4 <= {{(`LOG2_NBY2-6){1'b0}},{5{1'b1}},1'b0};            7  :  ohd6c4 <= {{(`LOG2_NBY2-7){1'b0}},{6{1'b1}},1'b0};            8  :  ohd6c4 <= {{(`LOG2_NBY2-8){1'b0}},{7{1'b1}},1'b0};            9  :  ohd6c4 <= {{(`LOG2_NBY2-9){1'b0}},{8{1'b1}},1'b0};            10 :  ohd6c4 <= {{(`LOG2_NBY2-10){1'b0}},{9{1'b1}},1'b0};            11 :  ohd6c4 <= {{(`LOG2_NBY2-11){1'b0}},{10{1'b1}},1'b0};            12 :  ohd6c4 <= {{(`LOG2_NBY2-12){1'b0}},{11{1'b1}},1'b0};            default : ohd6c4 <= `NUM_POINTS/2-2;         endcase      end
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            qi5137 <= 1'b0;            ip75347 <= 1'b0;         end else begin            qi5137 <= pf6b624==ohd6c4;            ip75347 <= an8511f==ohd6c4;         end      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)          pf6b624 <= {`LOG2_NBY2{1'b0}};         else if(qi5137)       pf6b624 <= {`LOG2_NBY2{1'b0}};         else if(xj50aed) pf6b624 <= pf6b624 + 1'b1;         else               pf6b624 <= {`LOG2_NBY2{1'b0}};      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn)       an8511f <= {`LOG2_NBY2{1'b0}};         else if(ip75347)    an8511f <= {`LOG2_NBY2{1'b0}};         else if(gda1ad8) an8511f <= an8511f + 1'b1;         else            an8511f <= {`LOG2_NBY2{1'b0}};      end
      ep2c58b_FFTC2048 ea62c5d(                     .rstn       (rstn       ),                     .clk        (clk        ),                     .din        (an8511f      ),                     .fn6e854     (fn6e854     ),                     .oh33d38      (uv54fa8     ),                     .dout       (hbd8934       )                  );
      tj389da_FFTC2048 cmc4ed7(                     .rstn       (rstn       ),                     .clk        (clk        ),                     .din        (pf6b624      ),                     .ld71789      (fn6e854     ),                     .dout       (qgc49a6    )                  );
`ifdef BIT_REVERSE
      tj389da_FFTC2048 en4ed13(                     .rstn       (rstn       ),                     .clk        (clk        ),                     .din        (an8511f      ),                     .ld71789      (fn6e854     ),                     .dout       (ym88a40    )                  );
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            for(en75165=0;en75165<`WR_LATENCY;en75165=en75165+1) aa31148[en75165] <= {`LOG2_NBY2{1'b0}};         else begin            aa31148[0] <= hbd8934;            for(en75165=1;en75165<`WR_LATENCY;en75165=en75165+1) aa31148[en75165] <= aa31148[en75165-1];         end      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) thf9dcf <= {`LOG2_NBY2{1'b0}};         else      thf9dcf <= ir26988 ? qgc49a6 : aa31148[`WR_LATENCY-1];      end
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            vv45201 <= 1'b0;            oh2900e <= 1'b0;         end else begin            vv45201 <= oh2900e;            oh2900e <= mt8576e;         end      end
`ifdef BIT_REVERSE
      always @(posedge clk or negedge rstn)      begin         if(!rstn)          cmcee7f <= {`LOG2_NBY2{1'b0}};         else if(vv45201) cmcee7f <= ym88a40;         else               cmcee7f <= hbd8934;      end
`else
      always @(posedge clk or negedge rstn)      begin         if(!rstn) cmcee7f <= {`LOG2_NBY2{1'b0}};         else      cmcee7f <= hbd8934;      end
`endif
`ifdef ADDRESS_OUT
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ld403aa[0] <= 1'b0;         else if(hbd8934=={ohd6c4[`LOG2_NBY2-1:1],1'b1} && oh2900e )            ld403aa[0] <= 1'b1;         else if(!oh2900e)            ld403aa[0] <= 1'b0;      end      always @(posedge clk or negedge rstn)      begin         if(!rstn) ld403aa[1] <= 7'h00;         else      ld403aa[1] <= ld403aa[0];      end      always @(posedge clk or negedge rstn)      begin         if(!rstn) for(en75165=0;en75165<7;en75165=en75165+1) ho48075[en75165] <= {`LOG2_N{1'b0}};         else begin            ho48075[0] <= ls1d56 & ykdbf27 & kq566a7 | gd9a9c1;            for(en75165=1;en75165<7;en75165=en75165+1) ho48075[en75165] <= ho48075[en75165-1];         end      end
`ifdef TRUNCATE
         assign oaddr = ho48075[4];
`else
         assign oaddr = ho48075[5];
`endif
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module tj389da_FFTC2048 (
                  rstn,                
                  clk,                 
                  din,                 
                  ld71789,               
                  dout                 
               );
input                   rstn;
input                   clk;
input [`LOG2_NBY2-1:0]  din;
input [3:0]             ld71789;
output[`LOG2_NBY2-1:0]  dout;
reg [`LOG2_NBY2-1:0]    dout;
wire[`LOG2_NBY2-1:0]    ui4cd61;
integer                 en75165;
assign ui4cd61 = din << ld71789;
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            dout <= {`LOG2_NBY2{1'b0}};         else            for(en75165=0;en75165<`LOG2_NBY2;en75165=en75165+1) dout[en75165] <= ui4cd61[`LOG2_NBY2-1-en75165];      end
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module ep2c58b_FFTC2048 (
                  rstn,             
                  clk,              
                  din,              
                  fn6e854,           
                  oh33d38,            
                  dout              
               ) ;
input                      rstn;
input                      clk;
input [`LOG2_NBY2-1:0]     din;
input [3:0]                fn6e854;
input [`STAGE_WIDTH-1:0]   oh33d38;
output[`LOG2_NBY2-1:0]     dout;
reg [`LOG2_NBY2-1:0]       dout;
reg [(2*`LOG2_NBY2)-1:0]   ui4cd61;
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
`ifdef NUM_POINTS_64
`endif
`ifdef NUM_POINTS_128
`endif
`ifdef NUM_POINTS_256
`endif
`ifdef NUM_POINTS_512
`endif
`ifdef NUM_POINTS_1024
`endif
`ifdef NUM_POINTS_2048
`endif
`ifdef NUM_POINTS_4096
`endif
`ifdef NUM_POINTS_8192
`endif
`ifdef NUM_POINTS_16384
`endif
      always @(posedge clk or negedge rstn)      begin         if(!rstn)            ui4cd61 <= 0;         else            ui4cd61 <= din << oh33d38;      end
`ifdef NUM_POINTS_64
      always @* dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];
`endif
`ifdef NUM_POINTS_128
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_256
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_512
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_1024
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            4  :  dout <= {4'h0,ui4cd61[`LOG2_NBY2-5:0]} | ui4cd61[(2*`LOG2_NBY2)-5:`LOG2_NBY2-4];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_2048
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            4  :  dout <= {4'h0,ui4cd61[`LOG2_NBY2-5:0]} | ui4cd61[(2*`LOG2_NBY2)-5:`LOG2_NBY2-4];            5  :  dout <= {5'h0,ui4cd61[`LOG2_NBY2-6:0]} | ui4cd61[(2*`LOG2_NBY2)-6:`LOG2_NBY2-5];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_4096
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            4  :  dout <= {4'h0,ui4cd61[`LOG2_NBY2-5:0]} | ui4cd61[(2*`LOG2_NBY2)-5:`LOG2_NBY2-4];            5  :  dout <= {5'h0,ui4cd61[`LOG2_NBY2-6:0]} | ui4cd61[(2*`LOG2_NBY2)-6:`LOG2_NBY2-5];            6  :  dout <= {6'h0,ui4cd61[`LOG2_NBY2-7:0]} | ui4cd61[(2*`LOG2_NBY2)-7:`LOG2_NBY2-6];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_8192
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            4  :  dout <= {4'h0,ui4cd61[`LOG2_NBY2-5:0]} | ui4cd61[(2*`LOG2_NBY2)-5:`LOG2_NBY2-4];            5  :  dout <= {5'h0,ui4cd61[`LOG2_NBY2-6:0]} | ui4cd61[(2*`LOG2_NBY2)-6:`LOG2_NBY2-5];            6  :  dout <= {6'h0,ui4cd61[`LOG2_NBY2-7:0]} | ui4cd61[(2*`LOG2_NBY2)-7:`LOG2_NBY2-6];            7  :  dout <= {7'h0,ui4cd61[`LOG2_NBY2-8:0]} | ui4cd61[(2*`LOG2_NBY2)-8:`LOG2_NBY2-7];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
`ifdef NUM_POINTS_16384
      always @*      begin         case(fn6e854)            0  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];            1  :  dout <= {1'b0,ui4cd61[`LOG2_NBY2-2:0]} | ui4cd61[(2*`LOG2_NBY2)-2:`LOG2_NBY2-1];            2  :  dout <= {2'h0,ui4cd61[`LOG2_NBY2-3:0]} | ui4cd61[(2*`LOG2_NBY2)-3:`LOG2_NBY2-2];            3  :  dout <= {3'h0,ui4cd61[`LOG2_NBY2-4:0]} | ui4cd61[(2*`LOG2_NBY2)-4:`LOG2_NBY2-3];            4  :  dout <= {4'h0,ui4cd61[`LOG2_NBY2-5:0]} | ui4cd61[(2*`LOG2_NBY2)-5:`LOG2_NBY2-4];            5  :  dout <= {5'h0,ui4cd61[`LOG2_NBY2-6:0]} | ui4cd61[(2*`LOG2_NBY2)-6:`LOG2_NBY2-5];            6  :  dout <= {6'h0,ui4cd61[`LOG2_NBY2-7:0]} | ui4cd61[(2*`LOG2_NBY2)-7:`LOG2_NBY2-6];            7  :  dout <= {7'h0,ui4cd61[`LOG2_NBY2-8:0]} | ui4cd61[(2*`LOG2_NBY2)-8:`LOG2_NBY2-7];            8  :  dout <= {8'h0,ui4cd61[`LOG2_NBY2-9:0]} | ui4cd61[(2*`LOG2_NBY2)-9:`LOG2_NBY2-8];            default  :  dout <= ui4cd61[`LOG2_NBY2-1:0] | ui4cd61[(2*`LOG2_NBY2)-1:`LOG2_NBY2];         endcase      end
`endif
   endmodule                                                                                       
`timescale 1 ns / 100 ps
module pu9646c_FFTC2048 (
               clk,                 
               rstn,                
               vka88c0,            
               ip44602,            
               thf9dcf,          
               cmcee7f,          
               db9e2c7,           
               lqf163e,           
               lf8b1f2,          
               tu58f97           
               );
input                         clk;
input                         rstn;
input                         vka88c0;
input                         ip44602;
input [`LOG2_N-2:0]           thf9dcf;
input [`LOG2_N-2:0]           cmcee7f;
input [`DATA_WIDTH2-1:0]      db9e2c7;
input [`DATA_WIDTH2-1:0]      lqf163e;
output[`DATA_WIDTH2-1:0]      lf8b1f2;
output[`DATA_WIDTH2-1:0]      tu58f97;
`ifdef USE_DIST_RAM
reg [`DATA_WIDTH2-1:0]        lf8b1f2;
reg [`DATA_WIDTH2-1:0]        tu58f97;
wire[`DATA_WIDTH2-1:0]        zm2a98f;
wire[`DATA_WIDTH2-1:0]        sh54c7b;
`else
wire[`DATA_WIDTH2-1:0]        lf8b1f2;
wire[`DATA_WIDTH2-1:0]        tu58f97;
`endif
`ifdef USE_DIST_RAM
`else
`endif
`ifdef USE_DIST_RAM
`else
`endif
            
`ifdef USE_DIST_RAM
      defparam gd8f701.pmi_addr_depth       = (`NUM_POINTS/2  );      defparam gd8f701.pmi_addr_width       = (`LOG2_N-1      );      defparam gd8f701.pmi_data_width       = `DATA_WIDTH2;      defparam gd8f701.pmi_regmode          = "reg";      defparam gd8f701.pmi_init_file        = "none";      defparam gd8f701.pmi_init_file_format = "binary";      defparam gd8f701.pmi_family           = `DEVICE_FAMILY;      defparam gd8f701.module_type          = "pmi_distributed_dpram";      pmi_distributed_dpram   gd8f701(                        .WrAddress  (thf9dcf ),                        .Data       (db9e2c7  ),                        .WrClock    (clk        ),                        .WE         (vka88c0   ),                        .WrClockEn  (1'b1       ),                        .RdAddress  (cmcee7f ),                        .RdClock    (clk        ),                        .RdClockEn  (1'b1       ),                        .Reset      (1'b0       ),                        .Q          (zm2a98f     )                     );
      defparam hq114b0.pmi_addr_depth       = (`NUM_POINTS/2  );      defparam hq114b0.pmi_addr_width       = (`LOG2_N-1      );      defparam hq114b0.pmi_data_width       = `DATA_WIDTH2;      defparam hq114b0.pmi_regmode          = "reg";      defparam hq114b0.pmi_init_file        = "none";      defparam hq114b0.pmi_init_file_format = "binary";      defparam hq114b0.pmi_family           = `DEVICE_FAMILY;      defparam hq114b0.module_type          = "pmi_distributed_dpram";      pmi_distributed_dpram   hq114b0(                        .WrAddress  (thf9dcf ),                        .Data       (lqf163e  ),                        .WrClock    (clk        ),                        .WE         (ip44602   ),                        .WrClockEn  (1'b1       ),                        .RdAddress  (cmcee7f ),                        .RdClock    (clk        ),                        .RdClockEn  (1'b1       ),                        .Reset      (1'b0       ),                        .Q          (sh54c7b     )                     );
      always @(posedge clk or negedge rstn)      begin         if(!rstn) begin            lf8b1f2 <= {`DATA_WIDTH2{1'b0}};            tu58f97 <= {`DATA_WIDTH2{1'b0}};         end else begin            lf8b1f2 <= zm2a98f;            tu58f97 <= sh54c7b;         end      end
`else
      defparam gd8f701.pmi_wr_addr_depth = (`NUM_POINTS/2);      defparam gd8f701.pmi_wr_addr_width = (`LOG2_N-1);      defparam gd8f701.pmi_wr_data_width = `DATA_WIDTH2;      defparam gd8f701.pmi_rd_addr_depth = (`NUM_POINTS/2);      defparam gd8f701.pmi_rd_addr_width = (`LOG2_N-1);      defparam gd8f701.pmi_rd_data_width = `DATA_WIDTH2;      defparam gd8f701.pmi_regmode = "reg";      defparam gd8f701.pmi_gsr = "disable";      defparam gd8f701.pmi_resetmode = "sync";      defparam gd8f701.pmi_family = `DEVICE_FAMILY;      defparam gd8f701.pmi_init_file = "none";      defparam gd8f701.pmi_init_file_format = "binary";      defparam gd8f701.module_type = "pmi_ram_dp";      pmi_ram_dp gd8f701(                        .Data       (db9e2c7  ),                        .WrAddress  (thf9dcf ),                        .RdAddress  (cmcee7f ),                        .WrClock    (clk        ),                        .RdClock    (clk        ),                        .WrClockEn  (1'b1       ),                        .RdClockEn  (1'b1       ),                        .WE         (vka88c0   ),                        .Reset      (1'b0       ),                        .Q          (lf8b1f2 )                     );
      defparam db3de49.pmi_wr_addr_depth = (`NUM_POINTS/2);      defparam db3de49.pmi_wr_addr_width = (`LOG2_N-1);      defparam db3de49.pmi_wr_data_width = `DATA_WIDTH2;      defparam db3de49.pmi_rd_addr_depth = (`NUM_POINTS/2);      defparam db3de49.pmi_rd_addr_width = (`LOG2_N-1);      defparam db3de49.pmi_rd_data_width = `DATA_WIDTH2;      defparam db3de49.pmi_regmode = "reg";      defparam db3de49.pmi_gsr = "disable";      defparam db3de49.pmi_resetmode = "sync";      defparam db3de49.pmi_family = `DEVICE_FAMILY;      defparam db3de49.pmi_init_file = "none";      defparam db3de49.pmi_init_file_format = "binary";      defparam db3de49.module_type = "pmi_ram_dp";      pmi_ram_dp db3de49(                        .Data       (lqf163e  ),                        .WrAddress  (thf9dcf ),                        .RdAddress  (cmcee7f ),                        .WrClock    (clk        ),                        .RdClock    (clk        ),                        .WrClockEn  (1'b1       ),                        .RdClockEn  (1'b1       ),                        .WE         (ip44602   ),                        .Reset      (1'b0       ),                        .Q          (tu58f97 )                     );
`endif
   endmodule                                                                                                   
`timescale 1 ns / 100 ps
module psdf6d3_FFTC2048 (
                  clk,               
                  rstn,              
               `ifdef DYNAMIC_POINTS
                  points,
                  pointset,
               `endif
               `ifdef MODE_PORT_READ
                  mode,              
                  modeset,           
               `endif
               `ifdef SFACT_PORT_READ
                  sfact,             
                  sfactset,          
               `endif
                  ibstart,           
                  dire,              
                  diim,              
   
               `ifdef BFPU_PRESENT
                  exponent,          
               `else
                  `ifdef SFACT_UNSCALE
                  `else
                     except,         
                  `endif
               `endif
                  rfib,              
                  ibend,             
                  obstart,           
                  outvalid,          
               `ifdef ADDRESS_OUT
                  oaddr,             
               `endif
                  dore,              
                  doim               
                 );
input                         clk;
input                         rstn;
`ifdef DYNAMIC_POINTS
input [`NFFT_WIDTH-1:0]       points;
input                         pointset;
`endif
`ifdef MODE_PORT_READ
input                         mode;
input                         modeset;
`endif
`ifdef SFACT_PORT_READ
input [`SFACT_WIDTH-1:0]      sfact;
input                         sfactset;
`endif
input                         ibstart;
input [`DIN_WIDTH-1:0]        dire;
input [`DIN_WIDTH-1:0]        diim;
`ifdef BFPU_PRESENT
output[`STAGE_WIDTH:0]        exponent;
`else
`ifdef SFACT_UNSCALE
`else
output                     except;
`endif
`endif
output                        rfib;
output                        ibend;
output                        obstart;
output                        outvalid;
`ifdef ADDRESS_OUT
output[`LOG2_N-1:0]           oaddr;
`endif
output[`DATA_WIDTH-1:0]       dore;
output[`DATA_WIDTH-1:0]       doim;
wire[`DIN_WIDTH-1:0]         co820d5;
wire[`DIN_WIDTH-1:0]         uk106a9;
`ifdef SFACT_PORT_READ
wire[`SFACT_WIDTH-1:0]        psca410;
wire                          th618fa;
`endif
`ifdef DYNAMIC_POINTS
wire[`NFFT_WIDTH-1:0]         fc15ca;
wire                          vi63eb6;
`endif
`ifdef MODE_PORT_READ
wire                          ne57290;
`endif
wire                          cb9041a;
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
wire[`DATA_WIDTH-1:0]   kd44c3b;
wire[`DATA_WIDTH-1:0]   do30eec;
wire[`DATA_WIDTH-1:0]   ec3bb19;
wire[`DATA_WIDTH-1:0]   zxec646;
wire                    jc52b77;
`ifdef FULL_WIDTH
`else
`endif
wire[`LOG2_NBY2-1:0]    tjb0a23;
wire[`STAGE_WIDTH-1:0]  uv54fa8;
`ifdef TMEM_ALL
wire[`LOG2_NBY2-1:0]    jc760c3;
`else
wire[`LOG2_NBY4-1:0]    jc760c3;
wire[`LOG2_NBY4-1:0]    lqeec18;
wire[1:0]               qi9dd83;
`endif
`ifdef TMEM_ALL
`else
`endif
wire[`TWID_WIDTH2-1:0]   hoc502a;
`ifdef TMEM_ALL
`else
`endif
wire[`DATA_WIDTH2-1:0]  hd28152;
wire[`DATA_WIDTH2-1:0]  fn40a97;
wire[`DATA_WIDTH-1:0]   go7788d;
wire[`DATA_WIDTH-1:0]   ukbc468;
wire[`DATA_WIDTH-1:0]   ipe2340;
wire[`DATA_WIDTH-1:0]   do11a04;
wire[`TWID_WIDTH-1:0]   jrbf099;
wire[`TWID_WIDTH-1:0]   czf84cf;
wire[`DATA_WIDTH+1:0]   vvc267c;
wire[`DATA_WIDTH+1:0]   tj133e7;
wire[`DATA_WIDTH+1:0]   fc99f3e;
wire[`DATA_WIDTH+1:0]   bycf9f2;
wire[`LOG2_N-6:0]          sw2bb74;
wire[1:0]                  aaacedc;
wire[`DATA_WIDTH+1:0]      gq3e49d;
wire[`DATA_WIDTH+1:0]      enf24e9;
wire[`DATA_WIDTH+1:0]      ie9274d;
wire[`DATA_WIDTH+1:0]      vk93a68;
wire[`LOG2_NBY2-1:0]       db288fc;
`ifdef BFPU_PRESENT
wire[`STAGE_WIDTH:0]       exponent;
`endif
`ifdef BIT_REVERSE
wire[`LOG2_NBY2-1:0]       an8511f;
`endif
wire                       uka9d85;
wire                       al4ec28;
wire                       fa76144;
wire                       qi1f9a5;
wire                       oh23014;
`ifdef BFPU_PRESENT
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`else
`endif
wire[`DATA_WIDTH-1:0]      zz91389;
wire[`DATA_WIDTH-1:0]      fc89c4f;
wire[`DATA_WIDTH-1:0]      yx4e27b;
wire[`DATA_WIDTH-1:0]      vv713dd;
wire                       vica285;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
wire[`DATA_WIDTH-1:0]      vv4f773;
wire[`DATA_WIDTH-1:0]      xj7bb9f;
wire[`DATA_WIDTH-1:0]      hbddcfe;
wire[`DATA_WIDTH-1:0]      rgee7f6;
wire                       uk3ea23;
wire                       pf742a7;
wire                       qva153e;
wire[`LOG2_NBY2-1:0]    thf9dcf;
wire[`LOG2_NBY2-1:0]    cmcee7f;
wire[`STAGE_WIDTH-1:0]  ne5dba1;
wire[`STAGE_WIDTH-1:0]  nga7d44;
wire[3:0]               fn6e854;
wire                    ir8a15d;
wire                    wj5142b;
wire                    xj50aed;
wire                    mt8576e;
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
wire[`DATA_WIDTH2-1:0]  cz6f567;
wire[`DATA_WIDTH2-1:0]  mr7ab3c;
wire[`DATA_WIDTH-1:0]      vid59e4;
wire[`DATA_WIDTH-1:0]      ukacf22;
wire                       gof5118;
`ifdef OUTVALID_SEL
`endif
wire                       ir95bbb;
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef FULL_WIDTH
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BIT_REVERSE
`endif
`ifdef BFPU_PRESENT
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`else
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef FULL_WIDTH
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef TMEM_ALL
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BIT_REVERSE
`endif
`ifdef BFPU_PRESENT
`ifdef BFPU_PRESENT
`ifdef BIT_REVERSE
`endif
`endif
`else
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BIT_REVERSE
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef OUTVALID_SEL
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`endif
`ifdef BFPU_PRESENT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef OUTVALID_SEL
`endif
      
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
         
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
         
`ifdef SFACT_PORT_READ
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
                  jpc7848_FFTC2048 vx2206b (                      .clk          (clk           ),                      .rstn         (rstn          ),
`ifdef DYNAMIC_POINTS
                      .points       (points        ),                      .xw48d1e   (pointset      ),
`endif
`ifdef MODE_PORT_READ
                      .mode         (mode          ),                      .co34798     (modeset       ),
`endif
`ifdef SFACT_PORT_READ
                      .sfact        (sfact         ),                      .do1e601    (sfactset      ),
`endif
                      .nrf300a     (ibstart       ),                      .co98057        (dire          ),                      .hoc02b9        (diim          ),
`ifdef DYNAMIC_POINTS
                      .fc15ca     (fc15ca      ),                      .ouae52 (vi63eb6   ),
`endif
`ifdef MODE_PORT_READ
                      .ne57290       (ne57290        ),                      .ieb9482   (ieb9482    ),
`endif
`ifdef SFACT_PORT_READ
                      .psca410      (psca410       ),                      .zk52083  (zk52083   ),
`endif
                      .cb9041a   (cb9041a    ),                      .co820d5      (co820d5       ),                      .uk106a9      (uk106a9       )                  );
         
`ifdef FULL_WIDTH
         assign kd44c3b = {{(`DATA_WIDTH-`DIN_WIDTH){co820d5[`DIN_WIDTH-1]}},co820d5};         assign do30eec = {{(`DATA_WIDTH-`DIN_WIDTH){uk106a9[`DIN_WIDTH-1]}},uk106a9};
`else
         assign kd44c3b = co820d5;         assign do30eec = uk106a9;
`endif
         sj12f6f_FFTC2048 rt6b283 (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .fft_mode      (jc52b77     ),                     .dire          (kd44c3b      ),                     .diim          (do30eec      ),                     .dore          (ec3bb19      ),                     .doim          (zxec646      )                 );
         
`ifdef TMEM_ALL
`else
`endif
         yx4b493_FFTC2048 bl7166f(                     .rstn          (rstn          ),                     .clk           (clk           ),                     .tjb0a23          (tjb0a23          ),                     .uv54fa8        (uv54fa8        ),
`ifdef TMEM_ALL
`else
                     .qi9dd83     (qi9dd83     ),                     .lqeec18        (lqeec18        ),
`endif
                     .jc760c3        (jc760c3        )                  ) ;
                  dmfb478_FFTC2048 suf55ba(                     .clk           (clk           ),                     .rstn          (rstn          ),                     .jc760c3        (jc760c3        ),
`ifdef TMEM_ALL
`else
                     .lqeec18        (lqeec18        ),                     .qi9dd83     (qi9dd83     ),
`endif
                     .aa1a145         (hoc502a         )                  );
                  assign jrbf099 = hoc502a[`TWID_WIDTH2-1:`TWID_WIDTH];         assign czf84cf = hoc502a[`TWID_WIDTH-1:0];         assign go7788d = hd28152[`DATA_WIDTH2-1:`DATA_WIDTH];         assign ukbc468 = hd28152[`DATA_WIDTH-1:0];         assign ipe2340 = fn40a97[`DATA_WIDTH2-1:`DATA_WIDTH];         assign do11a04 = fn40a97[`DATA_WIDTH-1:0];
         ec10059_FFTC2048 ohbbedd (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .pub262    (go7788d       ),                     .czc9899    (ukbc468       ),                     .yk59313    (ipe2340       ),                     .yk4c4cd    (do11a04       ),                     .os62668    (jrbf099       ),                     .bn13340    (czf84cf       ),                     .ri99a06   (vvc267c       ),                     .qg68196   (tj133e7       ),                     .vvcd032   (fc99f3e       ),                     .zx40cb1   (bycf9f2       )               ) ;
`ifdef BFPU_PRESENT
`endif
`ifdef BIT_REVERSE
`endif
`ifdef BFPU_PRESENT
         tw3016e_FFTC2048 en511d7 (                     .rstn          (rstn          ),                     .clk           (clk           ),                     .rv2dca9         (vvc267c       ),                     .dz6e54e         (tj133e7       ),                     .su72a76         (fc99f3e       ),                     .oh953b0         (bycf9f2       ),
`ifdef BFPU_PRESENT
                     .uka9d85  (uka9d85  ),                     .tjb0a23          (tjb0a23          ),
`ifdef BIT_REVERSE
                     .an8511f         (an8511f         ),
`endif
                     .db288fc        (db288fc        ),                     .al4ec28       (al4ec28       ),                     .fa76144       (fa76144       ),                     .exponent      (exponent      ),                     .cz709f8         (aaacedc        ),                     .qi1f9a5     (qi1f9a5     ),                     .ibend         (oh23014     ),                     .uv447e6        (uvd9450  ),
`endif
                     .ks34a7f         (gq3e49d     ),                     .hda53f9         (enf24e9     ),                     .an29fcf         (ie9274d     ),                     .xj4fe7c         (vk93a68     )                  );
`else
         assign gq3e49d = vvc267c;         assign enf24e9 = tj133e7;         assign ie9274d = fc99f3e;         assign vk93a68 = bycf9f2;
`endif
                  rtf9aaf_FFTC2048 nr610df (                     .rstn          (rstn          ),                     .clk           (clk           ),                     .cz709f8         (aaacedc        ),                     .vica285      (vica285      ),                     .rv2dca9         (gq3e49d     ),                     .dz6e54e         (enf24e9     ),                     .su72a76         (ie9274d     ),                     .oh953b0         (vk93a68     ),                     .go7788d       (go7788d       ),                     .ukbc468       (ukbc468       ),                     .ipe2340       (ipe2340       ),                     .do11a04       (do11a04       ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
                     .except        (dmfb548       ),
`endif
`endif
                     .ks34a7f         (zz91389      ),                     .hda53f9         (fc89c4f      ),                     .an29fcf         (yx4e27b      ),                     .xj4fe7c         (vv713dd      )                  );
                  sj232d3_FFTC2048 gbfdb8c (                     .rstn          (rstn          ),                     .clk           (clk           ),                     .uk3ea23          (uk3ea23          ),                     .end39ce     (ec3bb19      ),                     .tw9ce75     (zxec646      ),                     .rv2dca9         (zz91389      ),                     .dz6e54e         (fc89c4f      ),                     .su72a76         (yx4e27b      ),                     .oh953b0         (vv713dd      ),                     .pf742a7         (pf742a7         ),                     .qva153e         (qva153e         ),                     .ks34a7f         (vv4f773        ),                     .hda53f9         (xj7bb9f        ),                     .an29fcf         (hbddcfe        ),                     .xj4fe7c         (rgee7f6        )                  );
                  ba2adc0_FFTC2048 ri355cd (                     .rstn          (rstn          ),                     .clk           (clk           ),                     .ir8a15d       (ir8a15d       ),                     .wj5142b       (wj5142b       ),                     .xj50aed     (xj50aed     ),                     .mt8576e       (mt8576e       ),                     .fn6e854        (fn6e854        ),                     .uv54fa8        (uv54fa8        ),                     .ne5dba1      (ne5dba1      ),
`ifdef BIT_REVERSE
                     .an8511f         (an8511f         ),
`endif
`ifdef ADDRESS_OUT
                     .oaddr         (oaddr         ),
`endif
                     .thf9dcf    (thf9dcf    ),                     .cmcee7f    (cmcee7f    )                  );
                  assign cz6f567 = {vv4f773,xj7bb9f};         assign mr7ab3c = {hbddcfe,rgee7f6};         pu9646c_FFTC2048 zz69ac (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .vka88c0      (vka88c0      ),                     .ip44602      (ip44602      ),                     .thf9dcf    (thf9dcf    ),                     .cmcee7f    (cmcee7f    ),                     .db9e2c7     (cz6f567         ),                     .lqf163e     (mr7ab3c         ),                     .lf8b1f2    (hd28152        ),                     .tu58f97    (fn40a97        )                  );
                  epd4c0_FFTC2048 ieb6b7a (                     .rstn          (rstn          ),                     .clk           (clk           ),                     .aa98120           (gof5118          ),      
`ifdef OUTVALID_SEL
                     .ng14954        (ng14954        ),
`endif
                        .rv2dca9         (zz91389      ),                     .dz6e54e         (fc89c4f      ),                     .su72a76         (yx4e27b      ),                     .oh953b0         (vv713dd      ),                     .dore          (vid59e4      ),                     .doim          (ukacf22      )               );
                  sj12f6f_FFTC2048 ym92daa (                     .clk           (clk           ),                     .rstn          (rstn          ),                     .fft_mode      (ir95bbb     ),                     .dire          (vid59e4      ),                     .diim          (ukacf22      ),                     .dore          (dore          ),                     .doim          (doim          )                 );
                  ymb9ff3_FFTC2048 qi3e827 (                     .rstn          (rstn       ),                     .clk           (clk        ),                     .vife654   (cb9041a ),
`ifdef DYNAMIC_POINTS
                     .points        (fc15ca   ),                     .pu9951f     (vi63eb6),
`endif
`ifdef MODE_PORT_READ
                     .mode          (ne57290     ),                     .modeset       (ieb9482 ),
`endif
`ifdef SFACT_PORT_READ
                     .sfact         (psca410    ),                     .sfactset      (zk52083),
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
                     .dmfb548       (dmfb548    ),
`endif
`endif
                     .jc52b77     (jc52b77  ),                     .ir95bbb     (ir95bbb  ),
`ifdef BFPU_PRESENT
`else
                     .aaacedc        (aaacedc     ),
`endif
`ifdef BFPU_PRESENT
                     .al4ec28       (al4ec28    ),                     .fa76144       (fa76144    ),                     .uka9d85  (uka9d85  ),                     .qi1f9a5     (qi1f9a5  ),                     .uvd9450  (uvd9450),
`endif
                     .vica285      (vica285   ),                     .ir8a15d       (ir8a15d    ),                     .wj5142b       (wj5142b    ),                     .xj50aed     (xj50aed  ),                     .mt8576e       (mt8576e    ),                     .sw2bb74        (sw2bb74     ),                     .ne5dba1      (ne5dba1   ),                     .db288fc        (db288fc     ),                     .fn6e854        (fn6e854     ),                     .pf742a7         (pf742a7      ),                     .qva153e         (qva153e      ),                     .tjb0a23          (tjb0a23       ),                     .uv54fa8        (uv54fa8     ),                     .nga7d44        (nga7d44     ),                     .uk3ea23          (uk3ea23       ),                     .gof5118          (gof5118       ),                     .vka88c0      (vka88c0   ),                     .ip44602      (ip44602   ),                     .oh23014     (oh23014  ),
                     .rfib          (rfib       ),                     .ibend         (ibend      ),
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
                     .except        (except     ),
`endif
`endif
      
`ifdef OUTVALID_SEL
                     .ng14954        (ng14954     ),
`endif
                        .obstart       (obstart    ),                     .outvalid      (outvalid   )                  );
   endmodule
`endif
`timescale 1 ns / 100 ps
module FFTC2048 (
               clk,                 
               rstn,                
            `ifdef DYNAMIC_POINTS
               points,              
               pointset,            
            `endif
            `ifdef MODE_PORT_READ
               mode,                
               modeset,             
            `endif
            `ifdef SFACT_PORT_READ
               sfact,               
               sfactset,            
            `endif
               ibstart,             
               dire,                
               diim,                
            `ifdef BFPU_PRESENT
               exponent,            
            `else
               `ifdef SFACT_UNSCALE
               `else
                  except,              
               `endif
            `endif
               rfib,                
               ibend,               
               obstart,             
               outvalid,            
           `ifdef HP_FFT
           `else
                 `ifdef ADDRESS_OUT
                    oaddr,               
                 `endif
           `endif
                    dore,                
                    doim                 
                    )
   `ifdef DEVICE_ECP
    
   `else
   `ifdef DEVICE_ECP2
    
   `else
   `ifdef DEVICE_ECP3
    
   `else
   `ifdef DEVICE_ECP2M
    
   `else
   `ifdef DEVICE_XP2
    
   `else
    
   `endif
   `endif
   `endif
   `endif
   `endif
 ;
`ifdef HP_FFT
parameter pnfft_width  = `NFFT_WIDTH;
parameter pdin_widthr  = `DIN_WIDTH;
parameter ptwid_widthr = `TWID_WIDTH;
parameter pdout_widthr = `DOUT_WIDTH;
parameter pnum_points  = `NUM_POINTS;
parameter plog2_points = `LOG2_POINTS;
parameter fixed_scaling= `SCALE_VAL;
parameter device_family = `DEVICE_FAMILY;
`ifdef DYNAMIC_POINTS
parameter pdyn_points      = 1;
`else
parameter pdyn_points      = 0;
`endif
parameter sfact_width         = 2*plog2_points;
`ifdef TRUNCATE
parameter rounding_method  = 1;
`else
parameter rounding_method  = 0;
`endif
`ifdef BIT_REVERSE
parameter bit_reverse  = 1;
`else
parameter bit_reverse  = 0;
`endif
`ifdef MODE_FORWARD
parameter fft_mode     = 0;
`endif 
`ifdef MODE_INVERSE
parameter fft_mode     = 1;
`endif 
`ifdef MODE_PORT_READ
parameter fft_mode     = 2;
`endif 
`ifdef FULL_WAVE
parameter mem_type     = 0;
`endif 
`ifdef RQUARTER_WAVE
parameter mem_type     = 1;
`endif 
`ifdef CQUARTER_WAVE
parameter mem_type     = 2;
`endif 
`ifdef SUMOFANGLES_WAVE
parameter mem_type     = 3;
`endif 
`ifdef WMEM_DIST
parameter pebr_thresh = 9;
`endif
`ifdef WMEM_EBR
parameter pebr_thresh = 5;
`endif
`ifdef WMEM_AUTO
parameter pebr_thresh = 7;
`endif
`ifdef USE_HARDMAC
parameter phard_mac = 1;
`else
parameter phard_mac = 0;
`endif
`ifdef SCALE_REG
parameter pscale_reg = 1;
`else
parameter pscale_reg = 0;
`endif
`ifdef TRUNCATE_LASTSTGS
parameter ptrunc_laststgs = 1;
`else
parameter ptrunc_laststgs = 0;
`endif
`ifdef DYNAMIC_POINTS
parameter pbfimux_level   = `BFIMUX_LEVEL;
parameter pcntmux_level   = `CNTMUX_LEVEL;
`else
parameter pbfimux_level   = 0;
parameter pcntmux_level   = 0;
`endif
localparam co2b2ce      = 2*pdin_widthr;
localparam ng114ec     = 2*pdout_widthr;
localparam vve6110     = 2*ptwid_widthr;
localparam rtec748  = plog2_points-1;
input                                     clk;
input                                     rstn;
input                                     ibstart;
`ifdef DYNAMIC_POINTS
input [pnfft_width-1:0]                points;
input                                  pointset;
`endif
`ifdef MODE_PORT_READ
input                                  mode;
input                                  modeset;
`endif
`ifdef SFACT_PORT_READ
input [sfact_width-1:0]                sfact;
input                                  sfactset;
`endif
input  [pdin_widthr-1:0]                  dire;
input  [pdin_widthr-1:0]                  diim;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
output                              except;
`endif
`endif
output                                    ibend;
output                                    rfib;
output                                    outvalid;
output                                    obstart;
output [pdout_widthr-1:0]                 dore;
output [pdout_widthr-1:0]                 doim;
wire [sfact_width-1:0]                    vve93e5;
wire                                      kq49f2f;
wire [pnfft_width-1:0]                    fa7cbce;
wire                                      uie5e73;
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
wire                                except;
`endif
`endif
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef SFACT_PORT_READ
`else
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef MODE_FORWARD
`endif
`ifdef MODE_INVERSE
`endif
`else
input                      clk;
input                      rstn;
`ifdef DYNAMIC_POINTS
input [`NFFT_WIDTH-1:0]    points;
input                      pointset;
`endif
`ifdef MODE_PORT_READ
input                      mode;
input                      modeset;
`endif
`ifdef SFACT_PORT_READ
input [`SFACT_WIDTH-1:0]   sfact;
input                      sfactset;
`endif
input                      ibstart;
input [`DIN_WIDTH-1:0]     dire;
input [`DIN_WIDTH-1:0]     diim;
`ifdef BFPU_PRESENT
output[`STAGE_WIDTH:0]     exponent;
`else
`ifdef SFACT_UNSCALE
`else
output                  except;
`endif
`endif
output                     rfib;
output                     ibend;
output                     obstart;
output                     outvalid;
`ifdef ADDRESS_OUT
output[`LOG2_N-1:0]        oaddr;
`endif
output[`DATA_WIDTH-1:0]    dore;
output[`DATA_WIDTH-1:0]    doim;
`ifdef BFPU_PRESENT
wire[`STAGE_WIDTH:0]       exponent;
`else
`ifdef SFACT_UNSCALE
`else
wire                    except;
`endif
`endif
wire                       rfib;
wire                       ibend;
wire                       outvalid;
`ifdef ADDRESS_OUT
wire[`LOG2_N-1:0]          oaddr;
`endif
wire[`DATA_WIDTH-1:0]      dore;
wire[`DATA_WIDTH-1:0]      doim;
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`endif
`ifdef HP_FFT
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef MODE_FORWARD
`endif 
`ifdef MODE_INVERSE
`endif 
`ifdef MODE_PORT_READ
`endif 
`ifdef FULL_WAVE
`endif 
`ifdef RQUARTER_WAVE
`endif 
`ifdef CQUARTER_WAVE
`endif 
`ifdef SUMOFANGLES_WAVE
`endif 
`ifdef WMEM_DIST
`endif
`ifdef WMEM_EBR
`endif
`ifdef WMEM_AUTO
`endif
`ifdef USE_HARDMAC
`else
`endif
`ifdef SCALE_REG
`else
`endif
`ifdef TRUNCATE_LASTSTGS
`else
`endif
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef SFACT_PORT_READ
`else
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef MODE_FORWARD
`endif
`ifdef MODE_INVERSE
`endif
`else
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`endif
`ifdef HP_FFT
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef TRUNCATE
`else
`endif
`ifdef BIT_REVERSE
`else
`endif
`ifdef MODE_FORWARD
`endif 
`ifdef MODE_INVERSE
`endif 
`ifdef MODE_PORT_READ
`endif 
`ifdef FULL_WAVE
`endif 
`ifdef RQUARTER_WAVE
`endif 
`ifdef CQUARTER_WAVE
`endif 
`ifdef SUMOFANGLES_WAVE
`endif 
`ifdef WMEM_DIST
`endif
`ifdef WMEM_EBR
`endif
`ifdef WMEM_AUTO
`endif
`ifdef USE_HARDMAC
`else
`endif
`ifdef SCALE_REG
`else
`endif
`ifdef TRUNCATE_LASTSTGS
`else
`endif
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef DYNAMIC_POINTS
`else
`endif
`ifdef SFACT_PORT_READ
`else
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef MODE_FORWARD
`endif
`ifdef MODE_INVERSE
`endif
`else
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
`endif
`ifdef HP_FFT
                     
`ifdef DYNAMIC_POINTS
      
`else
      
`endif
   
`ifdef TRUNCATE
      
`else
      
`endif
`ifdef BIT_REVERSE
      
`else
      
`endif
`ifdef MODE_FORWARD
      
`endif 
`ifdef MODE_INVERSE
      
`endif 
`ifdef MODE_PORT_READ
      
`endif 
`ifdef FULL_WAVE
      
`endif 
`ifdef RQUARTER_WAVE
      
`endif 
`ifdef CQUARTER_WAVE
      
`endif 
`ifdef SUMOFANGLES_WAVE
      
`endif 
`ifdef WMEM_DIST
      
`endif
`ifdef WMEM_EBR
      
`endif
`ifdef WMEM_AUTO
      
`endif
`ifdef USE_HARDMAC
      
`else
      
`endif
`ifdef SCALE_REG
      
`else
      
`endif
`ifdef TRUNCATE_LASTSTGS
      
`else
      
`endif
`ifdef DYNAMIC_POINTS
            
`else
`endif
         
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
   
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
   
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef DYNAMIC_POINTS
      assign fa7cbce    = points;      assign uie5e73  = pointset;
`else
      assign fa7cbce    = 0;      assign uie5e73  = 1'b0;
`endif
`ifdef SFACT_PORT_READ
      assign vve93e5    = sfact;      assign kq49f2f = sfactset;
`else
      assign vve93e5    = 0;      assign kq49f2f = 1'b0;
`endif
`ifdef MODE_PORT_READ
      assign ymbc92f    = mode;      assign wy24bca = modeset;
`endif
`ifdef MODE_FORWARD
      assign ymbc92f    = 1'b0;      assign wy24bca = 1'b0;
`endif
`ifdef MODE_INVERSE
      assign ymbc92f    = 1'b1;      assign wy24bca = 1'b1;
`endif
      twbd919_FFTC2048 #(         .pnfft_width       (pnfft_width),         .pdyn_points       (pdyn_points),         .pdin_widthr       (pdin_widthr),         .ptwid_widthr      (ptwid_widthr),         .pdout_widthr      (pdout_widthr),         .pnum_points       (pnum_points),         .plog2_points      (plog2_points),         .fixed_scaling     (fixed_scaling),         .rounding_method   (rounding_method),         .device_family     (device_family),         .bit_reverse       (bit_reverse),         .fft_mode          (fft_mode),         .pfe3535         (mem_type),         .sfact_width       (sfact_width),         .pebr_thresh       (pebr_thresh),         .pscale_reg        (pscale_reg),         .ptrunc_laststgs   (ptrunc_laststgs),         .pbfimux_level     (pbfimux_level),         .pcntmux_level     (pcntmux_level),         .phard_mac         (phard_mac)         )        swa35b2 (         .clk               (clk),                  .rstn              (rstn),                 .ibstart           (ibstart),              .pointset          (uie5e73),            .points            (fa7cbce),              .modeset           (wy24bca),             .mode              (ymbc92f),                .sfact             (vve93e5),               .sfactset          (kq49f2f),            .dire              (dire),                 .diim              (diim),                 .ibend             (ibend),                .rfib              (rfib),                 .outvalid          (outvalid),             .obstart           (obstart),              .except            (except),               .dore              (dore),                 .doim              (doim)                  );
`else
      
`ifdef DYNAMIC_POINTS
`endif
`ifdef MODE_PORT_READ
`endif
`ifdef SFACT_PORT_READ
`endif
      
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
      
`ifdef BFPU_PRESENT
`else
`ifdef SFACT_UNSCALE
`else
`endif
`endif
`ifdef ADDRESS_OUT
`endif
      psdf6d3_FFTC2048 ng14bb7 (                      .clk                (clk        ),                      .rstn               (rstn       ),
`ifdef DYNAMIC_POINTS
                      .points             (points     ),                      .pointset           (pointset  ),
`endif
`ifdef MODE_PORT_READ
                      .mode               (mode       ),                      .modeset            (modeset    ),
`endif
`ifdef SFACT_PORT_READ
                      .sfact              (sfact      ),                      .sfactset           (sfactset   ),
`endif
                      .ibstart            (ibstart    ),                      .dire               (dire       ),                      .diim               (diim       ),
`ifdef BFPU_PRESENT
                      .exponent           (exponent   ),
`else
`ifdef SFACT_UNSCALE
`else
                         .except          (except     ),
`endif
`endif
                      .rfib               (rfib       ),                      .ibend              (ibend      ),                      .obstart            (obstart    ),                      .outvalid           (outvalid   ),
`ifdef ADDRESS_OUT
                      .oaddr              (oaddr      ),
`endif
                      .dore               (dore       ),                      .doim               (doim       )                    ) ;
`endif
endmodule
`timescale 1 ns / 100 ps
module descram_FFTC2048 ( din,  dout);
parameter SIZE = 2047;
parameter SCRAMSTRING = 0;
localparam [31:0] zkdfd9d = SCRAMSTRING;
localparam zxf675a = SCRAMSTRING & 4'hf;
localparam [11:0] co9d6b8 = 'h7ff;
input  [(1 << zxf675a)  -1:0] din;
output [SIZE-1:0] dout;
reg    [SIZE-1:0] dout;
reg [zxf675a-1:0] qvbe403 [0:1];
reg [zxf675a-1:0] an900ed;
reg oh8076d;
integer lf3b6c;
integer rtd7680;
   initial begin   lf3b6c = $fopen(".fred");   $fdisplay( lf3b6c, "%3h\n%3h", (zkdfd9d >> 4) & co9d6b8, (zkdfd9d >> (zxf675a+4)) & co9d6b8 );   $fclose(lf3b6c);   $readmemh(".fred", qvbe403);   end   always @ (din) begin   an900ed = qvbe403[1];       for (rtd7680=0; rtd7680<SIZE; rtd7680=rtd7680+1) begin           dout[rtd7680] = din[an900ed];       oh8076d  = ^(an900ed & qvbe403[0]);       an900ed =  {an900ed, oh8076d};       end   end endmodule
